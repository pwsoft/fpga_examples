library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

-- ------------------------------------------------------------------------

entity gigatron_tb_rom is
	port (
		a : in unsigned(15 downto 0);
		q : out unsigned(15 downto 0)
	);
end entity;

-- ------------------------------------------------------------------------

architecture rtl of gigatron_tb_rom is
	subtype rom_data_elem_t is unsigned(7 downto 0);
	type rom_data_t is array(integer range 0 to 65535) of rom_data_elem_t;
	signal rom_data_byte0 : rom_data_t := (
		X"00",X"18",X"18",X"C1",X"00",X"D6",X"00",X"69",
		X"CA",X"C2",X"69",X"EC",X"00",X"69",X"CA",X"61",
		X"F0",X"01",X"FC",X"82",X"00",X"C2",X"EC",X"A0",
		X"01",X"EC",X"A0",X"00",X"18",X"18",X"00",X"D2",
		X"D6",X"01",X"F4",X"8D",X"60",X"C2",X"01",X"F4",
		X"81",X"60",X"C2",X"81",X"C2",X"01",X"80",X"EC",
		X"D2",X"01",X"80",X"EC",X"D6",X"00",X"18",X"18",
		X"00",X"C2",X"90",X"00",X"D6",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"00",
		X"C2",X"00",X"C2",X"C2",X"C2",X"C2",X"C2",X"00",
		X"18",X"18",X"00",X"C2",X"C2",X"C2",X"00",X"18",
		X"18",X"C2",X"C2",X"14",X"E0",X"C2",X"00",X"C2",
		X"00",X"C2",X"14",X"CA",X"CA",X"CA",X"C2",X"C2",
		X"00",X"C2",X"00",X"C2",X"C2",X"C2",X"00",X"C2",
		X"00",X"C2",X"00",X"C2",X"01",X"A0",X"C2",X"14",
		X"E0",X"00",X"02",X"02",X"02",X"02",X"02",X"02",
		X"14",X"E0",X"00",X"14",X"E0",X"00",X"14",X"E0",
		X"00",X"14",X"E0",X"00",X"14",X"E0",X"00",X"14",
		X"E0",X"00",X"14",X"E0",X"00",X"14",X"E0",X"00",
		X"14",X"E0",X"00",X"14",X"E0",X"00",X"14",X"E0",
		X"00",X"14",X"E0",X"00",X"14",X"E0",X"00",X"14",
		X"E0",X"00",X"14",X"E0",X"00",X"14",X"E0",X"00",
		X"14",X"E0",X"00",X"14",X"E0",X"00",X"14",X"E0",
		X"00",X"14",X"E0",X"00",X"14",X"E0",X"00",X"14",
		X"E0",X"00",X"14",X"E0",X"00",X"14",X"E0",X"00",
		X"14",X"E0",X"00",X"14",X"E0",X"00",X"14",X"E0",
		X"00",X"14",X"E0",X"00",X"14",X"E0",X"00",X"14",
		X"E0",X"00",X"14",X"E0",X"00",X"14",X"E0",X"00",
		X"14",X"E0",X"00",X"14",X"E0",X"00",X"14",X"E0",
		X"00",X"14",X"E0",X"00",X"14",X"E0",X"15",X"14",
		X"E0",X"01",X"02",X"02",X"19",X"02",X"14",X"E0",
		X"00",X"C3",X"00",X"C2",X"02",X"14",X"E0",X"00",
		X"15",X"E0",X"00",X"00",X"C2",X"00",X"C2",X"00",
		X"C2",X"00",X"C2",X"81",X"C2",X"61",X"61",X"81",
		X"C2",X"81",X"C2",X"E8",X"FC",X"60",X"60",X"81",
		X"C2",X"01",X"F0",X"FC",X"A0",X"01",X"C2",X"F0",
		X"FC",X"00",X"00",X"81",X"EC",X"FC",X"00",X"E4",
		X"C2",X"80",X"FE",X"FC",X"00",X"C2",X"FC",X"21",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C2",X"00",X"C2",X"01",X"F0",X"00",X"C2",X"15",
		X"E0",X"00",X"14",X"E0",X"14",X"01",X"20",X"C2",
		X"01",X"EC",X"FC",X"00",X"00",X"41",X"C2",X"01",
		X"F0",X"FC",X"A0",X"00",X"C2",X"19",X"01",X"21",
		X"80",X"19",X"D6",X"00",X"29",X"89",X"CA",X"30",
		X"05",X"89",X"89",X"CA",X"20",X"69",X"12",X"09",
		X"14",X"8D",X"E8",X"FC",X"20",X"00",X"81",X"C2",
		X"01",X"14",X"19",X"01",X"F4",X"80",X"C2",X"A0",
		X"EC",X"A1",X"00",X"FC",X"C2",X"EC",X"00",X"FC",
		X"C2",X"01",X"02",X"60",X"C2",X"01",X"60",X"EC",
		X"FC",X"C3",X"C0",X"01",X"20",X"F0",X"01",X"00",
		X"C2",X"15",X"E0",X"00",X"FC",X"19",X"40",X"21",
		X"C2",X"C0",X"00",X"C2",X"15",X"E0",X"00",X"FC",
		X"19",X"E0",X"14",X"01",X"60",X"EC",X"01",X"A0",
		X"C2",X"20",X"F0",X"00",X"FC",X"FC",X"00",X"EC",
		X"A0",X"02",X"00",X"C2",X"FC",X"02",X"C2",X"00",
		X"C2",X"00",X"C2",X"01",X"60",X"EC",X"01",X"E8",
		X"01",X"C2",X"01",X"C2",X"FC",X"00",X"00",X"C2",
		X"C2",X"02",X"C2",X"00",X"EC",X"A0",X"02",X"C2",
		X"FC",X"00",X"01",X"20",X"C2",X"00",X"C2",X"15",
		X"E0",X"00",X"14",X"09",X"C2",X"C2",X"EC",X"FC",
		X"00",X"00",X"C2",X"01",X"21",X"80",X"14",X"E0",
		X"18",X"02",X"02",X"02",X"02",X"02",X"02",X"FC",
		X"01",X"00",X"C2",X"14",X"11",X"0D",X"DE",X"C2",
		X"0D",X"91",X"15",X"00",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"18",X"01",X"21",X"80",
		X"18",X"D6",X"00",X"29",X"89",X"CA",X"30",X"05",
		X"89",X"89",X"CA",X"20",X"69",X"12",X"09",X"14",
		X"8D",X"E8",X"FC",X"20",X"00",X"81",X"C2",X"01",
		X"FD",X"18",X"00",X"C2",X"14",X"01",X"90",X"01",
		X"8D",X"FD",X"D2",X"00",X"C2",X"01",X"40",X"21",
		X"C2",X"C0",X"FD",X"11",X"11",X"01",X"A0",X"F0",
		X"80",X"C2",X"00",X"FD",X"C2",X"C0",X"00",X"FD",
		X"C2",X"14",X"E0",X"00",X"01",X"80",X"D2",X"01",
		X"A5",X"F0",X"C2",X"FC",X"00",X"C2",X"00",X"C2",
		X"15",X"E0",X"00",X"02",X"02",X"02",X"02",X"FC",
		X"15",X"81",X"E8",X"C2",X"01",X"80",X"D2",X"0D",
		X"DE",X"FE",X"0D",X"80",X"E4",X"A0",X"14",X"E1",
		X"00",X"C2",X"DE",X"0D",X"C2",X"01",X"80",X"C2",
		X"00",X"FC",X"12",X"05",X"14",X"E0",X"C2",X"14",
		X"E0",X"12",X"80",X"C2",X"05",X"C2",X"11",X"05",
		X"C2",X"FC",X"00",X"12",X"80",X"C2",X"01",X"C6",
		X"11",X"01",X"C6",X"FC",X"00",X"01",X"EC",X"C2",
		X"01",X"F0",X"00",X"C2",X"0D",X"FE",X"01",X"EC",
		X"F0",X"0D",X"02",X"FC",X"0D",X"01",X"FC",X"80",
		X"DE",X"0D",X"C2",X"FC",X"00",X"F8",X"E4",X"0D",
		X"F4",X"E8",X"0D",X"E8",X"F4",X"0D",X"E4",X"F8",
		X"0D",X"C2",X"00",X"C2",X"FC",X"00",X"12",X"01",
		X"C6",X"FC",X"00",X"11",X"05",X"C2",X"01",X"90",
		X"05",X"C2",X"01",X"80",X"C2",X"01",X"A0",X"C2",
		X"FC",X"00",X"F0",X"EC",X"0D",X"01",X"B0",X"01",
		X"C6",X"01",X"A0",X"D2",X"01",X"FC",X"C6",X"15",
		X"E0",X"81",X"14",X"E0",X"21",X"14",X"E0",X"01",
		X"41",X"C2",X"FC",X"00",X"61",X"C2",X"FC",X"00",
		X"C2",X"FC",X"00",X"12",X"14",X"E0",X"00",X"14",
		X"E0",X"12",X"80",X"C2",X"01",X"85",X"C2",X"E8",
		X"A5",X"FC",X"45",X"25",X"02",X"30",X"05",X"81",
		X"11",X"85",X"C2",X"FC",X"00",X"14",X"E0",X"01",
		X"A0",X"C2",X"FC",X"00",X"81",X"E8",X"15",X"E1",
		X"12",X"80",X"C2",X"01",X"E8",X"A5",X"C2",X"FC",
		X"45",X"C2",X"25",X"02",X"30",X"01",X"A5",X"11",
		X"A5",X"C2",X"00",X"FC",X"15",X"14",X"E0",X"C2",
		X"01",X"80",X"C2",X"01",X"C2",X"11",X"05",X"A0",
		X"C2",X"01",X"90",X"05",X"D6",X"FC",X"00",X"81",
		X"C2",X"FC",X"00",X"14",X"E0",X"C2",X"14",X"E0",
		X"C2",X"14",X"E0",X"01",X"14",X"E0",X"14",X"E0",
		X"14",X"E0",X"C2",X"14",X"E0",X"C2",X"14",X"E0",
		X"14",X"E0",X"14",X"E0",X"14",X"E0",X"C2",X"01",
		X"A0",X"C2",X"01",X"C2",X"14",X"E0",X"00",X"01",
		X"80",X"C2",X"01",X"C2",X"01",X"C2",X"14",X"E0",
		X"00",X"02",X"C2",X"00",X"C2",X"14",X"E0",X"00",
		X"81",X"C2",X"E8",X"A1",X"FC",X"41",X"21",X"02",
		X"30",X"05",X"81",X"14",X"E0",X"C2",X"01",X"E8",
		X"A1",X"C2",X"FC",X"41",X"C2",X"21",X"02",X"30",
		X"01",X"A5",X"14",X"E0",X"C2",X"30",X"81",X"C2",
		X"05",X"81",X"81",X"C2",X"01",X"A0",X"14",X"E0",
		X"C2",X"81",X"C2",X"90",X"01",X"C6",X"11",X"01",
		X"C6",X"14",X"E0",X"00",X"81",X"C2",X"90",X"05",
		X"C2",X"11",X"05",X"C2",X"14",X"E0",X"00",X"90",
		X"05",X"16",X"11",X"05",X"12",X"01",X"CE",X"14",
		X"E0",X"00",X"A0",X"C2",X"11",X"15",X"0D",X"C2",
		X"00",X"C2",X"14",X"E0",X"00",X"90",X"05",X"16",
		X"11",X"05",X"12",X"01",X"DE",X"01",X"CE",X"14",
		X"E0",X"00",X"01",X"A0",X"C2",X"11",X"15",X"0D",
		X"DE",X"C2",X"0D",X"14",X"E0",X"C2",X"C2",X"90",
		X"05",X"21",X"C2",X"11",X"05",X"21",X"C2",X"14",
		X"E0",X"C2",X"90",X"05",X"41",X"C2",X"11",X"05",
		X"41",X"C2",X"14",X"E0",X"90",X"05",X"61",X"C2",
		X"11",X"05",X"61",X"C2",X"14",X"E0",X"00",X"01",
		X"61",X"61",X"81",X"C2",X"C2",X"81",X"C2",X"E8",
		X"FC",X"60",X"60",X"81",X"C2",X"C2",X"14",X"E0",
		X"00",X"01",X"30",X"01",X"82",X"45",X"C2",X"01",
		X"30",X"05",X"C2",X"14",X"E0",X"00",X"01",X"C2",
		X"00",X"C2",X"14",X"E0",X"00",X"01",X"C2",X"00",
		X"C2",X"14",X"E0",X"00",X"11",X"15",X"01",X"DE",
		X"01",X"DE",X"01",X"DE",X"01",X"DE",X"14",X"E0",
		X"00",X"14",X"E0",X"11",X"85",X"C6",X"14",X"E0",
		X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"01",X"C2",X"01",X"C2",X"01",X"C2",X"01",X"C2",
		X"14",X"E0",X"00",X"F0",X"90",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",
		X"02",X"14",X"00",X"C2",X"01",X"20",X"E2",X"FC",
		X"C2",X"01",X"20",X"80",X"20",X"41",X"C2",X"00",
		X"C2",X"01",X"20",X"E2",X"FC",X"C2",X"14",X"E0",
		X"00",X"14",X"00",X"C2",X"01",X"20",X"40",X"E2",
		X"FC",X"C2",X"01",X"82",X"82",X"82",X"82",X"82",
		X"82",X"41",X"C2",X"00",X"C2",X"01",X"20",X"40",
		X"E2",X"FC",X"C2",X"14",X"E0",X"00",X"14",X"00",
		X"C2",X"01",X"20",X"40",X"E2",X"FC",X"C2",X"01",
		X"82",X"82",X"82",X"82",X"82",X"41",X"C2",X"00",
		X"C2",X"01",X"20",X"40",X"E2",X"FC",X"C2",X"00",
		X"14",X"E0",X"14",X"00",X"C2",X"01",X"20",X"40",
		X"E2",X"FC",X"C2",X"01",X"82",X"82",X"82",X"82",
		X"41",X"C2",X"00",X"C2",X"01",X"20",X"40",X"E2",
		X"FC",X"C2",X"14",X"E0",X"00",X"14",X"00",X"C2",
		X"01",X"20",X"40",X"E2",X"FC",X"C2",X"01",X"82",
		X"82",X"82",X"41",X"C2",X"00",X"C2",X"01",X"20",
		X"40",X"E2",X"FC",X"C2",X"00",X"14",X"E0",X"14",
		X"00",X"C2",X"01",X"20",X"40",X"E2",X"FC",X"C2",
		X"01",X"82",X"82",X"41",X"C2",X"00",X"C2",X"01",
		X"20",X"40",X"E2",X"FC",X"C2",X"14",X"E0",X"00",
		X"14",X"00",X"C2",X"01",X"82",X"82",X"82",X"82",
		X"C2",X"01",X"20",X"40",X"E2",X"FC",X"41",X"C2",
		X"01",X"82",X"82",X"82",X"82",X"C2",X"00",X"14",
		X"E0",X"15",X"E0",X"01",X"C2",X"14",X"E0",X"00",
		X"14",X"01",X"50",X"0D",X"C2",X"01",X"20",X"82",
		X"82",X"82",X"82",X"C2",X"01",X"50",X"0D",X"50",
		X"0D",X"41",X"C2",X"01",X"20",X"82",X"82",X"C2",
		X"01",X"50",X"0D",X"50",X"0D",X"50",X"0D",X"41",
		X"C2",X"01",X"20",X"C2",X"14",X"E0",X"00",X"15",
		X"CE",X"C2",X"C2",X"14",X"00",X"E0",X"15",X"41",
		X"CE",X"C2",X"C2",X"14",X"E0",X"00",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"14",X"E0",X"01",X"01",X"FC",X"11",X"01",X"FC",
		X"60",X"14",X"E0",X"00",X"14",X"E0",X"00",X"14",
		X"E0",X"14",X"14",X"E0",X"14",X"14",X"E0",X"14",
		X"15",X"F8",X"A0",X"F4",X"C2",X"20",X"F0",X"01",
		X"DE",X"DE",X"DE",X"FC",X"DE",X"00",X"EC",X"A0",
		X"01",X"20",X"F0",X"01",X"DE",X"FC",X"DE",X"02",
		X"02",X"02",X"01",X"20",X"F0",X"FC",X"01",X"0D",
		X"CE",X"14",X"E0",X"00",X"02",X"C2",X"01",X"DE",
		X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"DE",X"01",
		X"80",X"C2",X"01",X"F0",X"FC",X"00",X"00",X"81",
		X"C2",X"14",X"E0",X"00",X"EC",X"FC",X"00",X"C2",
		X"01",X"F0",X"14",X"61",X"60",X"EC",X"FC",X"C2",
		X"02",X"E0",X"00",X"01",X"20",X"80",X"FE",X"FC",
		X"00",X"00",X"00",X"00",X"C2",X"01",X"20",X"80",
		X"FE",X"FC",X"00",X"00",X"00",X"00",X"C2",X"01",
		X"20",X"80",X"FE",X"FC",X"00",X"00",X"00",X"00",
		X"C2",X"E0",X"00",X"F0",X"11",X"01",X"A0",X"14",
		X"E0",X"C2",X"15",X"0D",X"21",X"EC",X"FC",X"00",
		X"00",X"C2",X"01",X"82",X"EC",X"FC",X"00",X"C2",
		X"20",X"81",X"D2",X"01",X"A0",X"F0",X"14",X"C2",
		X"01",X"60",X"F0",X"C2",X"C2",X"E0",X"00",X"01",
		X"A0",X"C2",X"E0",X"00",X"C2",X"C2",X"E0",X"00",
		X"80",X"C2",X"01",X"D6",X"0D",X"DE",X"A0",X"C2",
		X"0D",X"14",X"E0",X"C2",X"14",X"05",X"61",X"F4",
		X"01",X"E8",X"FC",X"00",X"00",X"85",X"C2",X"E0",
		X"14",X"05",X"61",X"F4",X"01",X"E8",X"FC",X"00",
		X"E0",X"00",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"11",X"15",X"0D",X"F4",X"DE",X"81",X"C2",X"01",
		X"80",X"C2",X"01",X"80",X"C2",X"02",X"14",X"E0",
		X"00",X"C2",X"0D",X"DE",X"C2",X"0D",X"DE",X"C2",
		X"0D",X"DE",X"C2",X"0D",X"DE",X"C2",X"0D",X"DE",
		X"C2",X"11",X"15",X"01",X"DE",X"01",X"DE",X"01",
		X"DE",X"01",X"DE",X"01",X"DE",X"01",X"DE",X"01",
		X"80",X"C2",X"01",X"80",X"C2",X"01",X"A0",X"C2",
		X"14",X"E0",X"00",X"02",X"02",X"02",X"02",X"02",
		X"11",X"15",X"0D",X"F4",X"DE",X"81",X"C2",X"01",
		X"A0",X"C2",X"01",X"80",X"C2",X"02",X"14",X"E0",
		X"00",X"C2",X"0D",X"DE",X"C2",X"0D",X"DE",X"C2",
		X"0D",X"DE",X"C2",X"0D",X"DE",X"C2",X"0D",X"DE",
		X"11",X"15",X"DE",X"01",X"DE",X"01",X"DE",X"01",
		X"DE",X"01",X"DE",X"01",X"DE",X"01",X"80",X"C2",
		X"01",X"80",X"C2",X"01",X"A0",X"C2",X"14",X"E0",
		X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"11",X"15",X"0D",X"F4",X"DE",X"60",X"80",X"81",
		X"C2",X"01",X"80",X"C2",X"01",X"80",X"C2",X"02",
		X"14",X"E0",X"00",X"C2",X"0D",X"DE",X"C2",X"0D",
		X"DE",X"C2",X"0D",X"DE",X"C2",X"0D",X"DE",X"C2",
		X"0D",X"DE",X"C2",X"11",X"15",X"01",X"DE",X"01",
		X"DE",X"01",X"DE",X"01",X"DE",X"01",X"DE",X"01",
		X"DE",X"01",X"80",X"C2",X"01",X"A0",X"C2",X"01",
		X"A0",X"C2",X"14",X"E0",X"00",X"02",X"02",X"02",
		X"11",X"15",X"0D",X"F4",X"DE",X"60",X"80",X"81",
		X"C2",X"01",X"A0",X"C2",X"01",X"80",X"C2",X"02",
		X"14",X"E0",X"00",X"C2",X"0D",X"DE",X"C2",X"0D",
		X"DE",X"C2",X"0D",X"DE",X"C2",X"0D",X"DE",X"C2",
		X"0D",X"DE",X"11",X"15",X"DE",X"01",X"DE",X"01",
		X"DE",X"01",X"DE",X"01",X"DE",X"01",X"DE",X"01",
		X"80",X"C2",X"01",X"A0",X"C2",X"01",X"A0",X"C2",
		X"14",X"E0",X"00",X"21",X"D2",X"14",X"CA",X"15",
		X"CD",X"01",X"EC",X"FC",X"01",X"C2",X"14",X"E0",
		X"00",X"09",X"C2",X"11",X"15",X"0D",X"D6",X"11",
		X"DD",X"DD",X"01",X"20",X"F0",X"FC",X"00",X"CD",
		X"81",X"81",X"D6",X"11",X"DD",X"DD",X"01",X"20",
		X"F0",X"FC",X"00",X"CD",X"81",X"81",X"D6",X"11",
		X"DD",X"DD",X"01",X"20",X"F0",X"FC",X"00",X"CD",
		X"81",X"81",X"D6",X"11",X"DD",X"DD",X"01",X"20",
		X"F0",X"FC",X"00",X"CD",X"81",X"81",X"D6",X"11",
		X"DD",X"DD",X"01",X"20",X"F0",X"FC",X"00",X"CD",
		X"81",X"81",X"D6",X"11",X"DD",X"DD",X"01",X"20",
		X"F0",X"FC",X"00",X"CD",X"81",X"81",X"D6",X"11",
		X"DD",X"DD",X"01",X"20",X"F0",X"FC",X"00",X"CD",
		X"81",X"81",X"D6",X"11",X"DD",X"DD",X"01",X"20",
		X"F0",X"FC",X"00",X"CD",X"81",X"81",X"11",X"15",
		X"CE",X"01",X"80",X"C2",X"61",X"F0",X"01",X"A0",
		X"C2",X"14",X"E0",X"00",X"14",X"E0",X"00",X"D6",
		X"00",X"E0",X"81",X"15",X"00",X"81",X"E8",X"01",
		X"20",X"80",X"20",X"C2",X"01",X"20",X"C2",X"0D",
		X"20",X"41",X"C2",X"00",X"C2",X"0D",X"20",X"14",
		X"E2",X"FC",X"14",X"E0",X"00",X"15",X"01",X"20",
		X"C2",X"0D",X"20",X"41",X"C2",X"00",X"C2",X"0D",
		X"20",X"14",X"E2",X"FC",X"15",X"0D",X"20",X"C2",
		X"01",X"20",X"8D",X"8D",X"CE",X"C2",X"C2",X"01",
		X"20",X"11",X"45",X"C2",X"14",X"00",X"E0",X"15",
		X"0D",X"20",X"C2",X"FC",X"00",X"02",X"01",X"C2",
		X"01",X"C2",X"14",X"E0",X"00",X"02",X"15",X"0D",
		X"DE",X"C2",X"0D",X"C2",X"14",X"E0",X"00",X"01",
		X"12",X"80",X"C2",X"05",X"C2",X"C2",X"C2",X"14",
		X"00",X"E0",X"14",X"01",X"A0",X"D2",X"01",X"C6",
		X"E0",X"00",X"00",X"C2",X"00",X"C2",X"14",X"00",
		X"E0",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"FC",
		X"A0",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"81",X"E8",X"C2",X"11",X"15",X"0D",X"C2",X"01",
		X"80",X"D2",X"F0",X"FC",X"00",X"00",X"81",X"D6",
		X"01",X"20",X"FE",X"FC",X"0D",X"01",X"E8",X"01",
		X"FC",X"00",X"80",X"E4",X"A0",X"00",X"C2",X"14",
		X"E1",X"00",X"02",X"02",X"01",X"C2",X"01",X"D2",
		X"80",X"C2",X"F0",X"FC",X"00",X"00",X"81",X"C2",
		X"FC",X"00",X"00",X"D2",X"00",X"C2",X"00",X"FC",
		X"02",X"FC",X"00",X"FC",X"81",X"FC",X"02",X"D2",
		X"00",X"C2",X"00",X"81",X"C2",X"F0",X"FC",X"00",
		X"00",X"81",X"C2",X"FC",X"00",X"F0",X"FC",X"00",
		X"00",X"81",X"C2",X"01",X"A0",X"C2",X"FC",X"00",
		X"FC",X"00",X"FC",X"01",X"01",X"C2",X"00",X"81",
		X"E8",X"01",X"01",X"60",X"F0",X"FC",X"01",X"01",
		X"8D",X"C2",X"E8",X"AD",X"FC",X"4D",X"2D",X"02",
		X"30",X"05",X"C2",X"01",X"80",X"D2",X"F0",X"FC",
		X"00",X"00",X"81",X"D6",X"0D",X"81",X"C2",X"01",
		X"80",X"C2",X"F0",X"FC",X"00",X"00",X"81",X"C2",
		X"11",X"FC",X"00",X"12",X"14",X"00",X"81",X"02",
		X"E8",X"01",X"80",X"C2",X"F0",X"FC",X"00",X"00",
		X"81",X"C2",X"0D",X"DE",X"C2",X"0D",X"C2",X"01",
		X"81",X"C2",X"E8",X"A1",X"FC",X"41",X"21",X"02",
		X"30",X"05",X"81",X"C2",X"11",X"FC",X"00",X"D2",
		X"E8",X"FC",X"00",X"00",X"C2",X"01",X"80",X"C2",
		X"F0",X"FC",X"00",X"00",X"81",X"C2",X"FC",X"00",
		X"81",X"C2",X"90",X"05",X"C2",X"11",X"05",X"D2",
		X"01",X"80",X"C2",X"F0",X"FC",X"00",X"00",X"81",
		X"C2",X"00",X"81",X"E8",X"C2",X"14",X"E1",X"FC",
		X"80",X"E4",X"A0",X"00",X"C2",X"14",X"E1",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",
		X"14",X"15",X"21",X"81",X"F0",X"8D",X"C2",X"C2",
		X"61",X"C2",X"0D",X"61",X"21",X"20",X"C2",X"01",
		X"C2",X"E8",X"AD",X"FC",X"4D",X"2D",X"02",X"30",
		X"01",X"20",X"45",X"41",X"C2",X"14",X"E0",X"00",
		X"C2",X"C2",X"C2",X"01",X"20",X"C2",X"14",X"00",
		X"E0",X"15",X"0D",X"60",X"C2",X"00",X"D2",X"00",
		X"C2",X"00",X"C2",X"14",X"E0",X"00",X"01",X"FC",
		X"20",X"01",X"40",X"C2",X"02",X"E0",X"00",X"01",
		X"E8",X"F4",X"01",X"F4",X"E8",X"01",X"20",X"F0",
		X"EC",X"01",X"20",X"EC",X"F0",X"01",X"20",X"F0",
		X"EC",X"01",X"20",X"EC",X"F0",X"01",X"F0",X"EC",
		X"01",X"EC",X"F0",X"01",X"81",X"C2",X"E8",X"A1",
		X"FC",X"41",X"21",X"02",X"30",X"05",X"81",X"81",
		X"C2",X"02",X"E0",X"00",X"02",X"01",X"80",X"C2",
		X"C2",X"C2",X"00",X"E0",X"02",X"E0",X"00",X"01",
		X"A0",X"FC",X"C2",X"01",X"80",X"FC",X"C2",X"01",
		X"A0",X"FC",X"C2",X"00",X"E0",X"15",X"01",X"FC",
		X"2D",X"15",X"01",X"FC",X"4D",X"15",X"01",X"6D",
		X"C2",X"C2",X"C2",X"14",X"00",X"E0",X"14",X"E0",
		X"14",X"E0",X"01",X"A0",X"D2",X"14",X"01",X"C2",
		X"01",X"C2",X"80",X"C2",X"DE",X"F0",X"FC",X"00",
		X"00",X"81",X"C2",X"CE",X"11",X"15",X"0D",X"11",
		X"C2",X"15",X"0D",X"C2",X"14",X"00",X"E0",X"14",
		X"E0",X"14",X"E0",X"14",X"E0",X"14",X"E0",X"14",
		X"E0",X"14",X"E0",X"14",X"E0",X"14",X"E0",X"14",
		X"E0",X"14",X"E0",X"14",X"E0",X"14",X"E0",X"14",
		X"E0",X"14",X"E0",X"14",X"E0",X"14",X"E0",X"14",
		X"E0",X"14",X"E0",X"14",X"E0",X"14",X"E0",X"14",
		X"E0",X"14",X"E0",X"14",X"E0",X"14",X"E0",X"14",
		X"E0",X"14",X"E0",X"14",X"E0",X"14",X"E0",X"14",
		X"E0",X"14",X"E0",X"14",X"E0",X"14",X"E0",X"14",
		X"E0",X"14",X"E0",X"14",X"E0",X"14",X"E0",X"A0",
		X"C2",X"11",X"14",X"E1",X"FC",X"15",X"0D",X"A0",
		X"CE",X"C2",X"C2",X"14",X"00",X"E0",X"15",X"0D",
		X"80",X"CE",X"C2",X"C2",X"14",X"00",X"E0",X"02",
		X"02",X"15",X"0D",X"C2",X"C2",X"C2",X"02",X"14",
		X"E0",X"00",X"15",X"0D",X"FC",X"C2",X"15",X"0D",
		X"FC",X"C2",X"01",X"A1",X"91",X"05",X"C2",X"C2",
		X"C2",X"14",X"E0",X"00",X"15",X"01",X"CE",X"14",
		X"E0",X"00",X"15",X"01",X"CE",X"14",X"E0",X"00",
		X"01",X"A1",X"91",X"01",X"C6",X"14",X"E0",X"00",
		X"15",X"01",X"CE",X"14",X"E0",X"00",X"01",X"C2",
		X"C2",X"C2",X"14",X"E0",X"00",X"01",X"A0",X"C2",
		X"C2",X"C2",X"02",X"14",X"E0",X"00",X"01",X"80",
		X"FC",X"C2",X"01",X"FC",X"C2",X"01",X"FC",X"C2",
		X"01",X"FC",X"C2",X"01",X"FC",X"20",X"01",X"FC",
		X"40",X"01",X"FC",X"20",X"01",X"FC",X"40",X"01",
		X"20",X"C2",X"14",X"00",X"E0",X"02",X"11",X"15",
		X"0D",X"C2",X"21",X"C2",X"01",X"20",X"C2",X"0D",
		X"82",X"20",X"41",X"C2",X"14",X"E0",X"00",X"01",
		X"12",X"80",X"C2",X"14",X"0D",X"DE",X"80",X"C2",
		X"F0",X"FC",X"00",X"00",X"8D",X"C2",X"02",X"14",
		X"E0",X"00",X"01",X"A0",X"D2",X"01",X"20",X"F4",
		X"FC",X"60",X"C6",X"01",X"F0",X"FC",X"00",X"00",
		X"45",X"C6",X"01",X"20",X"45",X"40",X"C6",X"02",
		X"14",X"E0",X"00",X"FC",X"01",X"FC",X"01",X"01",
		X"15",X"E8",X"AD",X"C2",X"C2",X"FC",X"4D",X"C2",
		X"C2",X"2D",X"02",X"60",X"30",X"01",X"20",X"45",
		X"C2",X"14",X"E0",X"00",X"01",X"12",X"80",X"C2",
		X"05",X"C2",X"20",X"60",X"C2",X"05",X"20",X"80",
		X"C2",X"14",X"E0",X"00",X"01",X"12",X"80",X"C2",
		X"05",X"C2",X"20",X"60",X"C2",X"14",X"0D",X"DE",
		X"20",X"80",X"C2",X"0D",X"DE",X"C2",X"0D",X"C2",
		X"02",X"14",X"E0",X"00",X"02",X"02",X"02",X"02",
		X"09",X"49",X"EC",X"01",X"00",X"C2",X"15",X"E0",
		X"00",X"C2",X"01",X"C2",X"01",X"C2",X"01",X"C2",
		X"09",X"A0",X"C2",X"09",X"C2",X"01",X"C2",X"00",
		X"C2",X"00",X"C2",X"00",X"C2",X"15",X"E0",X"00",
		X"05",X"C2",X"01",X"C2",X"01",X"C2",X"01",X"C2",
		X"01",X"C2",X"02",X"14",X"E0",X"01",X"01",X"80",
		X"21",X"EC",X"01",X"80",X"21",X"EC",X"00",X"02",
		X"FC",X"A1",X"21",X"C2",X"01",X"41",X"C2",X"01",
		X"E0",X"C2",X"00",X"61",X"41",X"21",X"41",X"02",
		X"02",X"FC",X"02",X"D6",X"01",X"A0",X"D2",X"80",
		X"C2",X"DC",X"DC",X"80",X"DE",X"DC",X"DC",X"DC",
		X"DE",X"DC",X"DC",X"DC",X"DE",X"DC",X"DC",X"DC",
		X"DE",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"DC",X"80",X"DE",X"DC",X"80",X"DE",
		X"DC",X"DC",X"80",X"DE",X"DC",X"DC",X"80",X"DE",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"80",
		X"DE",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"DC",X"DC",X"14",X"E0",X"00",X"00",
		X"C2",X"95",X"01",X"E8",X"FC",X"01",X"01",X"CE",
		X"01",X"82",X"C2",X"01",X"81",X"94",X"01",X"E8",
		X"FC",X"01",X"01",X"CE",X"01",X"82",X"C2",X"01",
		X"A0",X"EC",X"80",X"14",X"E0",X"00",X"01",X"82",
		X"92",X"01",X"DE",X"20",X"EC",X"01",X"FC",X"81",
		X"60",X"DE",X"01",X"20",X"EC",X"FC",X"00",X"00",
		X"DE",X"01",X"CE",X"80",X"C2",X"60",X"F0",X"FC",
		X"00",X"00",X"81",X"C2",X"14",X"E0",X"00",X"11",
		X"0D",X"C2",X"11",X"0D",X"11",X"CE",X"82",X"82",
		X"81",X"C2",X"11",X"01",X"CE",X"01",X"80",X"C2",
		X"F0",X"FC",X"00",X"00",X"81",X"C2",X"14",X"E0",
		X"00",X"00",X"C2",X"01",X"D2",X"0D",X"C2",X"01",
		X"80",X"D2",X"0D",X"11",X"C6",X"01",X"80",X"C2",
		X"01",X"EC",X"A0",X"02",X"02",X"02",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"00",X"C2",X"00",X"14",X"E0",X"C2",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"15",X"0D",X"C2",X"A1",X"11",X"15",X"CE",
		X"01",X"A0",X"C2",X"01",X"C2",X"01",X"80",X"C2",
		X"EC",X"01",X"FC",X"02",X"A0",X"C2",X"14",X"E0",
		X"00",X"01",X"20",X"EC",X"FC",X"00",X"00",X"C2",
		X"15",X"01",X"80",X"D2",X"60",X"C2",X"C2",X"01",
		X"20",X"81",X"CE",X"01",X"80",X"C2",X"14",X"E0",
		X"00",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"00",X"C2",X"00",X"14",X"E0",X"C2",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"DC",X"00",X"C2",X"00",X"14",X"E0",
		X"C2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"00",X"C2",X"00",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"61",X"EC",X"11",X"15",X"03",X"CE",X"81",X"C2",
		X"01",X"80",X"C2",X"14",X"E0",X"00",X"01",X"A0",
		X"C2",X"14",X"E0",X"00",X"15",X"01",X"EC",X"01",
		X"B0",X"0D",X"DE",X"60",X"EC",X"0D",X"DE",X"20",
		X"C2",X"8D",X"80",X"20",X"C2",X"0D",X"DE",X"C2",
		X"0D",X"DE",X"C2",X"A0",X"20",X"41",X"EC",X"FC",
		X"00",X"00",X"21",X"C2",X"01",X"EC",X"01",X"C2",
		X"A0",X"C2",X"01",X"C2",X"C2",X"14",X"E0",X"00",
		X"00",X"EC",X"A0",X"02",X"00",X"C2",X"14",X"E0",
		X"00",X"01",X"B0",X"0D",X"C2",X"14",X"E0",X"00",
		X"01",X"F0",X"A0",X"C2",X"11",X"15",X"0D",X"11",
		X"15",X"CE",X"01",X"80",X"C2",X"FC",X"14",X"00",
		X"EC",X"A0",X"E0",X"00",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"DC",X"DC",X"00",X"C2",X"00",X"14",
		X"E0",X"C2",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"00",X"C2",X"00",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"DC",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"00",X"C2",
		X"00",X"14",X"E0",X"C2",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"00",X"C2",X"00",
		X"14",X"E0",X"C2",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"00",X"C2",X"00",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"DC",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"00",X"C2",
		X"00",X"14",X"E0",X"C2",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"DC",X"00",X"C2",X"00",X"14",X"E0",
		X"C2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"00",X"C2",X"00",X"14",X"E0",X"C2",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"00",X"C2",X"00",X"14",X"E0",X"C2",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"DC",X"00",X"C2",X"00",X"14",X"E0",
		X"C2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"00",
		X"C2",X"00",X"14",X"E0",X"C2",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"DC",X"DC",X"DC",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"00",X"C2",X"00",
		X"14",X"E0",X"C2",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"DC",X"00",X"C2",X"00",X"14",X"E0",X"C2",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"02",X"FE",X"FC",X"14",X"E0",X"C2",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"00",X"C2",X"00",X"14",X"E0",X"C2",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"FC",X"14",X"E0",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"10",X"16",
		X"01",X"A0",X"E2",X"14",X"00",X"14",X"E2",X"14",
		X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",
		X"00",X"C2",X"00",X"14",X"E0",X"C2",X"14",X"E0",
		X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"FE",X"FC",X"14",X"E0",X"C2",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		others => (others => '0'));
	signal rom_data_byte1 : rom_data_t := (
		X"00",X"80",X"C0",X"7C",X"01",X"01",X"FF",X"00",
		X"00",X"00",X"00",X"0B",X"FF",X"00",X"00",X"00",
		X"14",X"01",X"05",X"00",X"FF",X"00",X"16",X"01",
		X"00",X"15",X"01",X"01",X"80",X"C0",X"00",X"18",
		X"19",X"06",X"25",X"00",X"BF",X"06",X"07",X"2A",
		X"06",X"C1",X"07",X"08",X"08",X"18",X"01",X"21",
		X"18",X"19",X"01",X"21",X"19",X"03",X"80",X"C0",
		X"EE",X"16",X"02",X"01",X"17",X"59",X"5E",X"2B",
		X"22",X"B4",X"E2",X"00",X"00",X"FC",X"00",X"02",
		X"05",X"FF",X"0E",X"0F",X"10",X"11",X"12",X"07",
		X"80",X"C0",X"00",X"00",X"02",X"2C",X"0F",X"80",
		X"C0",X"13",X"14",X"01",X"03",X"2E",X"40",X"21",
		X"00",X"1C",X"01",X"F9",X"F6",X"F7",X"2C",X"1A",
		X"02",X"1B",X"F6",X"0A",X"0B",X"0C",X"AD",X"22",
		X"0E",X"24",X"F9",X"25",X"16",X"02",X"16",X"03",
		X"00",X"EA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"CB",X"F6",X"03",X"CB",X"F6",X"03",X"CB",
		X"F6",X"03",X"CB",X"F6",X"03",X"CB",X"F6",X"03",
		X"CB",X"F6",X"03",X"CB",X"F6",X"03",X"CB",X"F6",
		X"03",X"CB",X"F6",X"03",X"CB",X"F6",X"03",X"CB",
		X"F6",X"03",X"CB",X"F6",X"03",X"CB",X"F6",X"03",
		X"CB",X"F6",X"03",X"CB",X"F6",X"12",X"4B",X"00",
		X"03",X"CB",X"F6",X"03",X"CB",X"F6",X"03",X"CB",
		X"F6",X"03",X"CB",X"F6",X"03",X"CB",X"F6",X"03",
		X"CB",X"F6",X"03",X"CB",X"F6",X"03",X"CB",X"F6",
		X"03",X"CB",X"F6",X"03",X"CB",X"F6",X"03",X"CB",
		X"F6",X"03",X"CB",X"F6",X"03",X"CB",X"F6",X"03",
		X"CB",X"F6",X"03",X"CB",X"F6",X"03",X"CB",X"F6",
		X"03",X"CB",X"F6",X"03",X"CB",X"F6",X"03",X"CB",
		X"F6",X"03",X"CB",X"F6",X"12",X"E9",X"1B",X"FB",
		X"D5",X"19",X"00",X"00",X"24",X"00",X"03",X"CB",
		X"F5",X"18",X"00",X"19",X"00",X"03",X"CB",X"F4",
		X"05",X"FF",X"7F",X"C0",X"1F",X"80",X"20",X"B3",
		X"09",X"01",X"80",X"0E",X"0E",X"07",X"0F",X"06",
		X"06",X"08",X"08",X"16",X"17",X"53",X"6C",X"07",
		X"07",X"2D",X"1D",X"1E",X"01",X"2F",X"2D",X"22",
		X"23",X"00",X"01",X"2E",X"27",X"28",X"E8",X"2C",
		X"2E",X"48",X"00",X"48",X"0F",X"2E",X"48",X"14",
		X"0F",X"07",X"03",X"01",X"02",X"04",X"08",X"04",
		X"02",X"01",X"03",X"07",X"0F",X"0E",X"0C",X"08",
		X"04",X"02",X"01",X"02",X"04",X"08",X"0C",X"0E",
		X"14",X"10",X"0D",X"0E",X"52",X"55",X"1E",X"05",
		X"FF",X"23",X"12",X"00",X"01",X"21",X"FB",X"21",
		X"2C",X"5C",X"5D",X"00",X"F0",X"14",X"14",X"2C",
		X"63",X"64",X"01",X"00",X"2C",X"1F",X"02",X"21",
		X"01",X"20",X"02",X"7F",X"FE",X"FC",X"FE",X"80",
		X"00",X"FF",X"FD",X"FF",X"FC",X"FB",X"00",X"FA",
		X"07",X"00",X"7D",X"7E",X"3F",X"3F",X"03",X"03",
		X"13",X"12",X"1F",X"09",X"B1",X"02",X"09",X"BD",
		X"8D",X"0D",X"40",X"92",X"1F",X"91",X"C0",X"93",
		X"1F",X"1F",X"00",X"40",X"20",X"09",X"CF",X"9A",
		X"9B",X"0F",X"00",X"09",X"06",X"A6",X"03",X"A4",
		X"1E",X"05",X"FF",X"35",X"66",X"1F",X"0F",X"14",
		X"13",X"03",X"AF",X"1E",X"05",X"FF",X"33",X"66",
		X"1F",X"2E",X"01",X"11",X"EF",X"BE",X"12",X"01",
		X"12",X"7F",X"C6",X"EE",X"C5",X"C4",X"01",X"BF",
		X"01",X"00",X"80",X"12",X"CB",X"00",X"16",X"01",
		X"17",X"02",X"05",X"11",X"DF",X"E2",X"0B",X"D5",
		X"0A",X"0B",X"0C",X"0A",X"DA",X"F6",X"0A",X"0B",
		X"0A",X"00",X"0C",X"35",X"DC",X"01",X"00",X"11",
		X"EA",X"00",X"02",X"03",X"02",X"EA",X"1E",X"05",
		X"FF",X"26",X"01",X"F9",X"09",X"1F",X"F1",X"F2",
		X"01",X"EC",X"0D",X"02",X"21",X"01",X"02",X"B1",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"AE",
		X"02",X"CA",X"0D",X"01",X"09",X"00",X"00",X"20",
		X"00",X"1F",X"20",X"C0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"02",X"21",X"01",
		X"80",X"02",X"7F",X"FE",X"FC",X"FE",X"80",X"00",
		X"FF",X"FD",X"FF",X"FC",X"FB",X"00",X"FA",X"07",
		X"00",X"C4",X"C5",X"3F",X"3F",X"03",X"03",X"13",
		X"0D",X"C0",X"D3",X"0D",X"01",X"09",X"01",X"1F",
		X"00",X"0A",X"1F",X"DC",X"0D",X"03",X"0F",X"14",
		X"13",X"03",X"0B",X"1F",X"1F",X"09",X"EE",X"E5",
		X"F0",X"09",X"01",X"0C",X"0D",X"03",X"E9",X"0C",
		X"0D",X"01",X"04",X"C0",X"20",X"80",X"20",X"1F",
		X"00",X"F4",X"1F",X"F6",X"01",X"0D",X"FF",X"1E",
		X"05",X"FF",X"3C",X"00",X"00",X"00",X"00",X"03",
		X"17",X"15",X"0B",X"15",X"16",X"02",X"16",X"00",
		X"00",X"00",X"00",X"0E",X"0C",X"01",X"01",X"1E",
		X"00",X"18",X"00",X"00",X"19",X"16",X"01",X"16",
		X"F6",X"01",X"00",X"00",X"04",X"13",X"18",X"0B",
		X"BC",X"00",X"01",X"1D",X"00",X"18",X"1D",X"00",
		X"19",X"01",X"F6",X"00",X"01",X"1D",X"18",X"00",
		X"1D",X"19",X"00",X"01",X"F6",X"19",X"40",X"1D",
		X"18",X"43",X"01",X"1D",X"00",X"00",X"1D",X"45",
		X"48",X"00",X"00",X"3D",X"00",X"16",X"4A",X"01",
		X"00",X"00",X"16",X"01",X"F2",X"45",X"48",X"00",
		X"45",X"48",X"00",X"45",X"48",X"00",X"45",X"48",
		X"00",X"18",X"00",X"19",X"00",X"F8",X"00",X"18",
		X"00",X"00",X"F8",X"1C",X"00",X"1A",X"1C",X"01",
		X"00",X"1B",X"1C",X"02",X"1C",X"16",X"01",X"16",
		X"00",X"F3",X"45",X"48",X"00",X"1C",X"01",X"1B",
		X"00",X"1C",X"02",X"1C",X"1A",X"6D",X"00",X"19",
		X"FB",X"18",X"04",X"11",X"18",X"0B",X"B0",X"16",
		X"18",X"18",X"01",X"F9",X"18",X"18",X"01",X"F9",
		X"16",X"00",X"F9",X"00",X"04",X"E4",X"01",X"0B",
		X"C8",X"00",X"01",X"1D",X"18",X"00",X"18",X"A3",
		X"00",X"A5",X"00",X"00",X"00",X"80",X"00",X"19",
		X"1D",X"00",X"19",X"01",X"F2",X"04",X"62",X"16",
		X"02",X"16",X"CB",X"F6",X"15",X"AF",X"23",X"22",
		X"00",X"01",X"1D",X"18",X"C1",X"00",X"18",X"C4",
		X"00",X"18",X"00",X"00",X"80",X"19",X"00",X"1D",
		X"00",X"19",X"F2",X"01",X"17",X"04",X"07",X"1D",
		X"16",X"02",X"1A",X"17",X"1B",X"1D",X"00",X"02",
		X"16",X"1D",X"01",X"00",X"17",X"01",X"F3",X"1C",
		X"1C",X"01",X"F9",X"04",X"18",X"1D",X"04",X"26",
		X"1D",X"04",X"35",X"18",X"04",X"41",X"04",X"4C",
		X"04",X"57",X"1D",X"04",X"6D",X"1D",X"04",X"7A",
		X"04",X"86",X"04",X"91",X"04",X"9C",X"1D",X"1A",
		X"02",X"16",X"1B",X"17",X"03",X"CB",X"F6",X"16",
		X"02",X"18",X"17",X"19",X"1D",X"16",X"03",X"00",
		X"F4",X"00",X"18",X"00",X"19",X"03",X"CB",X"F5",
		X"18",X"18",X"1E",X"1D",X"20",X"1D",X"1D",X"00",
		X"80",X"00",X"19",X"03",X"CA",X"19",X"18",X"2C",
		X"1D",X"18",X"2F",X"1D",X"18",X"1D",X"00",X"80",
		X"19",X"00",X"03",X"CA",X"19",X"80",X"18",X"18",
		X"00",X"19",X"19",X"19",X"16",X"01",X"03",X"CA",
		X"16",X"1C",X"1D",X"01",X"19",X"00",X"1D",X"18",
		X"00",X"03",X"CB",X"F3",X"1C",X"1D",X"01",X"00",
		X"19",X"1D",X"00",X"18",X"03",X"CB",X"F3",X"01",
		X"00",X"00",X"1D",X"00",X"00",X"18",X"00",X"03",
		X"CB",X"F3",X"01",X"16",X"18",X"19",X"00",X"18",
		X"00",X"19",X"03",X"CB",X"F3",X"01",X"00",X"00",
		X"1D",X"00",X"00",X"18",X"00",X"19",X"00",X"03",
		X"CB",X"F2",X"16",X"01",X"16",X"18",X"19",X"00",
		X"00",X"18",X"00",X"03",X"CA",X"19",X"1D",X"01",
		X"00",X"19",X"19",X"1D",X"00",X"18",X"18",X"03",
		X"CA",X"1D",X"01",X"00",X"19",X"19",X"1D",X"00",
		X"18",X"18",X"03",X"CA",X"01",X"00",X"19",X"19",
		X"1D",X"00",X"18",X"18",X"03",X"CB",X"F3",X"0E",
		X"07",X"0F",X"06",X"06",X"18",X"08",X"08",X"B2",
		X"B3",X"53",X"6C",X"07",X"07",X"19",X"03",X"CB",
		X"EF",X"18",X"80",X"19",X"00",X"00",X"18",X"19",
		X"80",X"00",X"19",X"03",X"CB",X"F1",X"19",X"18",
		X"00",X"19",X"03",X"CB",X"F4",X"18",X"19",X"00",
		X"18",X"03",X"CB",X"F4",X"28",X"29",X"24",X"00",
		X"25",X"00",X"26",X"00",X"27",X"00",X"03",X"CB",
		X"F1",X"12",X"8F",X"28",X"00",X"00",X"03",X"00",
		X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"16",X"31",X"17",X"32",X"18",X"33",X"19",
		X"03",X"CB",X"F2",X"F0",X"01",X"12",X"20",X"1D",
		X"00",X"00",X"01",X"00",X"02",X"01",X"03",X"00",
		X"04",X"02",X"05",X"01",X"06",X"03",X"07",X"00",
		X"08",X"04",X"09",X"02",X"0A",X"05",X"0B",X"01",
		X"0C",X"06",X"0D",X"03",X"0E",X"07",X"0F",X"00",
		X"10",X"08",X"11",X"04",X"12",X"09",X"13",X"02",
		X"14",X"0A",X"15",X"05",X"16",X"0B",X"17",X"01",
		X"18",X"0C",X"19",X"06",X"1A",X"0D",X"1B",X"03",
		X"1C",X"0E",X"1D",X"07",X"1E",X"0F",X"1F",X"00",
		X"20",X"10",X"21",X"08",X"22",X"11",X"23",X"04",
		X"24",X"12",X"25",X"09",X"26",X"13",X"27",X"02",
		X"28",X"14",X"29",X"0A",X"2A",X"15",X"2B",X"05",
		X"2C",X"16",X"2D",X"0B",X"2E",X"17",X"2F",X"01",
		X"30",X"18",X"31",X"0C",X"32",X"19",X"33",X"06",
		X"34",X"1A",X"35",X"0D",X"36",X"1B",X"37",X"03",
		X"38",X"1C",X"39",X"0E",X"3A",X"1D",X"3B",X"07",
		X"3C",X"1E",X"3D",X"0F",X"3E",X"1F",X"3F",X"01",
		X"40",X"20",X"41",X"10",X"42",X"21",X"43",X"08",
		X"44",X"22",X"45",X"11",X"46",X"23",X"47",X"04",
		X"48",X"24",X"49",X"12",X"4A",X"25",X"4B",X"09",
		X"4C",X"26",X"4D",X"13",X"4E",X"27",X"4F",X"02",
		X"50",X"28",X"51",X"14",X"52",X"29",X"53",X"0A",
		X"54",X"2A",X"55",X"15",X"56",X"2B",X"57",X"05",
		X"58",X"2C",X"59",X"16",X"5A",X"2D",X"5B",X"0B",
		X"5C",X"2E",X"5D",X"17",X"5E",X"2F",X"5F",X"02",
		X"60",X"30",X"61",X"18",X"62",X"31",X"63",X"0C",
		X"64",X"32",X"65",X"19",X"66",X"33",X"67",X"06",
		X"68",X"34",X"69",X"1A",X"6A",X"35",X"6B",X"0D",
		X"6C",X"36",X"6D",X"1B",X"6E",X"37",X"6F",X"03",
		X"70",X"38",X"71",X"1C",X"72",X"39",X"73",X"0E",
		X"74",X"3A",X"75",X"1D",X"76",X"3B",X"77",X"07",
		X"78",X"3C",X"79",X"1E",X"7A",X"3D",X"7B",X"0F",
		X"7C",X"3E",X"7D",X"1F",X"7E",X"3F",X"7F",X"1D",
		X"00",X"05",X"08",X"1D",X"18",X"FE",X"00",X"FF",
		X"18",X"19",X"01",X"7F",X"80",X"18",X"18",X"15",
		X"1D",X"19",X"FE",X"00",X"FF",X"19",X"03",X"CB",
		X"E8",X"05",X"21",X"1D",X"18",X"FC",X"01",X"00",
		X"FF",X"18",X"19",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"18",X"32",X"1D",X"19",X"FC",X"01",
		X"00",X"FF",X"19",X"03",X"CB",X"E6",X"05",X"3E",
		X"1D",X"18",X"F8",X"03",X"00",X"FF",X"18",X"19",
		X"00",X"00",X"00",X"00",X"00",X"18",X"18",X"4E",
		X"1D",X"19",X"F8",X"03",X"00",X"FF",X"19",X"E6",
		X"03",X"CB",X"05",X"5A",X"1D",X"18",X"F0",X"07",
		X"00",X"FF",X"18",X"19",X"00",X"00",X"00",X"00",
		X"18",X"18",X"69",X"1D",X"19",X"F0",X"07",X"00",
		X"FF",X"19",X"03",X"CB",X"E7",X"05",X"75",X"1D",
		X"18",X"E0",X"0F",X"00",X"FF",X"18",X"19",X"00",
		X"00",X"00",X"18",X"18",X"83",X"1D",X"19",X"E0",
		X"0F",X"00",X"FF",X"19",X"E7",X"03",X"CB",X"05",
		X"8F",X"1D",X"18",X"C0",X"1F",X"00",X"FF",X"18",
		X"19",X"00",X"00",X"18",X"18",X"9C",X"1D",X"19",
		X"C0",X"1F",X"00",X"FF",X"19",X"03",X"CB",X"E8",
		X"05",X"AE",X"1D",X"19",X"00",X"00",X"00",X"00",
		X"19",X"18",X"F0",X"07",X"00",X"FF",X"19",X"19",
		X"18",X"00",X"00",X"00",X"00",X"18",X"E9",X"03",
		X"CB",X"2B",X"79",X"2A",X"26",X"03",X"CB",X"EC",
		X"07",X"26",X"03",X"00",X"27",X"26",X"03",X"00",
		X"00",X"00",X"00",X"26",X"25",X"03",X"00",X"03",
		X"00",X"26",X"26",X"25",X"0F",X"00",X"00",X"25",
		X"24",X"03",X"00",X"03",X"00",X"03",X"00",X"25",
		X"25",X"24",X"3F",X"24",X"03",X"CB",X"E4",X"25",
		X"00",X"28",X"29",X"0E",X"ED",X"20",X"25",X"19",
		X"00",X"28",X"29",X"0E",X"20",X"E9",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",
		X"00",X"00",X"A0",X"C0",X"00",X"A0",X"C0",X"28",
		X"FE",X"28",X"FE",X"28",X"24",X"54",X"FE",X"54",
		X"48",X"C4",X"C8",X"10",X"26",X"46",X"6C",X"92",
		X"6A",X"04",X"0A",X"00",X"A0",X"C0",X"00",X"00",
		X"00",X"38",X"44",X"82",X"00",X"00",X"82",X"44",
		X"38",X"00",X"28",X"10",X"7C",X"10",X"28",X"10",
		X"10",X"7C",X"10",X"10",X"00",X"05",X"06",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"02",
		X"02",X"00",X"00",X"00",X"06",X"18",X"60",X"00",
		X"7C",X"8A",X"92",X"A2",X"7C",X"22",X"42",X"FE",
		X"02",X"02",X"46",X"8A",X"92",X"92",X"62",X"44",
		X"82",X"92",X"92",X"6C",X"18",X"28",X"48",X"FE",
		X"08",X"E4",X"A2",X"A2",X"A2",X"9C",X"3C",X"52",
		X"92",X"92",X"0C",X"80",X"8E",X"90",X"A0",X"C0",
		X"6C",X"92",X"92",X"92",X"6C",X"60",X"92",X"92",
		X"94",X"78",X"00",X"24",X"24",X"00",X"00",X"00",
		X"25",X"26",X"00",X"00",X"10",X"28",X"44",X"82",
		X"00",X"28",X"28",X"28",X"28",X"28",X"00",X"82",
		X"44",X"28",X"10",X"40",X"80",X"8A",X"90",X"60",
		X"7C",X"82",X"BA",X"AA",X"78",X"3E",X"48",X"88",
		X"48",X"3E",X"FE",X"92",X"92",X"92",X"6C",X"7C",
		X"82",X"82",X"82",X"44",X"FE",X"82",X"82",X"44",
		X"38",X"FE",X"92",X"92",X"92",X"82",X"FE",X"90",
		X"90",X"90",X"80",X"7C",X"82",X"82",X"92",X"5C",
		X"FE",X"10",X"10",X"10",X"FE",X"00",X"82",X"FE",
		X"82",X"00",X"04",X"02",X"82",X"FC",X"80",X"FE",
		X"10",X"28",X"44",X"82",X"FE",X"02",X"02",X"02",
		X"02",X"FE",X"40",X"30",X"40",X"FE",X"FE",X"20",
		X"10",X"08",X"FE",X"7C",X"82",X"82",X"82",X"7C",
		X"FE",X"90",X"90",X"90",X"60",X"7C",X"82",X"8A",
		X"84",X"7A",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"FE",X"90",X"98",X"94",X"62",X"62",X"92",X"92",
		X"92",X"0C",X"80",X"80",X"FE",X"80",X"80",X"FC",
		X"02",X"02",X"02",X"FC",X"F0",X"0C",X"02",X"0C",
		X"F0",X"FE",X"04",X"18",X"04",X"FE",X"C6",X"28",
		X"10",X"28",X"C6",X"E0",X"10",X"0E",X"10",X"E0",
		X"86",X"8A",X"92",X"A2",X"C2",X"00",X"FE",X"82",
		X"82",X"00",X"00",X"60",X"18",X"06",X"00",X"00",
		X"82",X"82",X"FE",X"00",X"20",X"40",X"80",X"40",
		X"20",X"02",X"02",X"02",X"02",X"02",X"00",X"00",
		X"C0",X"A0",X"00",X"04",X"2A",X"2A",X"2A",X"1E",
		X"FE",X"22",X"22",X"22",X"1C",X"1C",X"22",X"22",
		X"22",X"02",X"1C",X"22",X"22",X"22",X"FE",X"1C",
		X"2A",X"2A",X"2A",X"18",X"10",X"7E",X"90",X"80",
		X"40",X"18",X"25",X"25",X"25",X"1E",X"FE",X"20",
		X"20",X"20",X"1E",X"00",X"22",X"BE",X"02",X"00",
		X"02",X"01",X"21",X"BE",X"00",X"FE",X"08",X"18",
		X"24",X"02",X"00",X"82",X"FE",X"02",X"00",X"3E",
		X"20",X"1C",X"20",X"1E",X"3E",X"10",X"20",X"20",
		X"1E",X"1C",X"22",X"22",X"22",X"1C",X"3F",X"24",
		X"24",X"24",X"18",X"18",X"24",X"24",X"24",X"3F",
		X"3E",X"10",X"20",X"20",X"10",X"12",X"2A",X"2A",
		X"2A",X"04",X"20",X"FC",X"22",X"02",X"04",X"3C",
		X"02",X"02",X"04",X"3E",X"38",X"04",X"02",X"04",
		X"38",X"3C",X"02",X"0C",X"02",X"3C",X"22",X"14",
		X"08",X"14",X"22",X"38",X"05",X"05",X"05",X"3E",
		X"22",X"26",X"2A",X"32",X"22",X"10",X"6C",X"82",
		X"82",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",
		X"82",X"82",X"6C",X"10",X"40",X"80",X"40",X"20",
		X"40",X"FE",X"FE",X"FE",X"FE",X"FE",X"10",X"38",
		X"54",X"10",X"10",X"10",X"20",X"7C",X"20",X"10",
		X"10",X"10",X"54",X"38",X"10",X"10",X"08",X"7C",
		X"08",X"10",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"00",X"00",X"45",X"00",X"49",X"00",X"4D",X"00",
		X"52",X"00",X"56",X"00",X"5C",X"00",X"61",X"00",
		X"67",X"00",X"6D",X"00",X"73",X"00",X"7A",X"00",
		X"01",X"01",X"09",X"01",X"11",X"01",X"1A",X"01",
		X"23",X"01",X"2D",X"01",X"37",X"01",X"42",X"01",
		X"4E",X"01",X"5A",X"01",X"67",X"01",X"74",X"01",
		X"03",X"02",X"12",X"02",X"23",X"02",X"34",X"02",
		X"46",X"02",X"5A",X"02",X"6E",X"02",X"04",X"03",
		X"1B",X"03",X"33",X"03",X"4D",X"03",X"69",X"03",
		X"06",X"04",X"25",X"04",X"45",X"04",X"68",X"04",
		X"0C",X"05",X"33",X"05",X"5C",X"05",X"08",X"06",
		X"36",X"06",X"67",X"06",X"1B",X"07",X"52",X"07",
		X"0C",X"08",X"49",X"08",X"0B",X"09",X"50",X"09",
		X"19",X"0A",X"67",X"0A",X"39",X"0B",X"10",X"0C",
		X"6C",X"0C",X"4E",X"0D",X"35",X"0E",X"23",X"0F",
		X"17",X"10",X"13",X"11",X"15",X"12",X"1F",X"13",
		X"32",X"14",X"4D",X"15",X"72",X"16",X"20",X"18",
		X"58",X"19",X"1C",X"1B",X"6B",X"1C",X"46",X"1E",
		X"2F",X"20",X"25",X"22",X"2A",X"24",X"3F",X"26",
		X"64",X"28",X"1A",X"2B",X"63",X"2D",X"3F",X"30",
		X"31",X"33",X"38",X"36",X"56",X"39",X"0D",X"3D",
		X"5E",X"40",X"4B",X"44",X"55",X"48",X"7E",X"4C",
		X"48",X"51",X"34",X"56",X"46",X"5B",X"7F",X"60",
		X"61",X"66",X"6F",X"6C",X"2C",X"73",X"1A",X"7A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"FF",X"EF",X"E2",X"D6",X"CB",X"C2",X"B9",X"B1",
		X"A9",X"A2",X"9C",X"96",X"91",X"8C",X"87",X"83",
		X"7F",X"7B",X"77",X"74",X"70",X"6D",X"6A",X"68",
		X"65",X"62",X"60",X"5E",X"5C",X"5A",X"58",X"56",
		X"54",X"52",X"50",X"4F",X"4D",X"4C",X"4A",X"49",
		X"48",X"46",X"45",X"44",X"43",X"42",X"41",X"40",
		X"3F",X"3E",X"3D",X"3C",X"3B",X"3A",X"39",X"38",
		X"37",X"37",X"36",X"35",X"34",X"34",X"33",X"32",
		X"32",X"31",X"30",X"30",X"2F",X"2F",X"2E",X"2E",
		X"2D",X"2D",X"2C",X"2C",X"2B",X"2B",X"2A",X"2A",
		X"29",X"29",X"28",X"28",X"27",X"27",X"27",X"26",
		X"26",X"26",X"25",X"25",X"24",X"24",X"24",X"23",
		X"23",X"23",X"22",X"22",X"22",X"22",X"21",X"21",
		X"21",X"20",X"20",X"20",X"20",X"1F",X"1F",X"1F",
		X"1F",X"1E",X"1E",X"1E",X"1E",X"1D",X"1D",X"1D",
		X"1D",X"1C",X"1C",X"1C",X"1C",X"1C",X"1B",X"1B",
		X"1B",X"1B",X"1B",X"1A",X"1A",X"1A",X"1A",X"1A",
		X"19",X"19",X"19",X"19",X"19",X"19",X"18",X"18",
		X"18",X"18",X"18",X"18",X"17",X"17",X"17",X"17",
		X"17",X"17",X"17",X"16",X"16",X"16",X"16",X"16",
		X"16",X"16",X"16",X"15",X"15",X"15",X"15",X"15",
		X"15",X"15",X"15",X"14",X"14",X"14",X"14",X"14",
		X"14",X"14",X"14",X"14",X"13",X"13",X"13",X"13",
		X"13",X"13",X"13",X"13",X"13",X"12",X"12",X"12",
		X"12",X"12",X"12",X"12",X"12",X"12",X"12",X"12",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"00",X"FD",X"04",X"68",X"18",
		X"0B",X"54",X"1E",X"24",X"18",X"26",X"09",X"83",
		X"B3",X"0C",X"FB",X"FC",X"0D",X"7F",X"0D",X"12",
		X"AE",X"07",X"12",X"CF",X"07",X"0D",X"09",X"01",
		X"27",X"3C",X"08",X"3E",X"24",X"04",X"25",X"25",
		X"00",X"00",X"00",X"28",X"00",X"01",X"26",X"01",
		X"24",X"02",X"2F",X"25",X"00",X"32",X"00",X"00",
		X"00",X"00",X"24",X"01",X"37",X"38",X"25",X"00",
		X"00",X"03",X"00",X"E8",X"00",X"24",X"25",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"26",
		X"08",X"26",X"24",X"4E",X"4F",X"FE",X"00",X"16",
		X"16",X"03",X"CB",X"E9",X"57",X"57",X"03",X"1E",
		X"19",X"63",X"03",X"18",X"B0",X"60",X"61",X"1E",
		X"00",X"CB",X"EF",X"18",X"03",X"68",X"00",X"6C",
		X"0A",X"0A",X"F6",X"F6",X"0A",X"18",X"03",X"72",
		X"00",X"76",X"0A",X"0A",X"0A",X"F6",X"0B",X"18",
		X"03",X"7C",X"00",X"80",X"0A",X"F6",X"F6",X"F6",
		X"0C",X"CB",X"E7",X"8A",X"24",X"16",X"02",X"03",
		X"CA",X"16",X"25",X"00",X"26",X"90",X"91",X"0E",
		X"12",X"0D",X"26",X"00",X"97",X"97",X"01",X"26",
		X"01",X"24",X"24",X"27",X"01",X"AC",X"03",X"27",
		X"0F",X"FF",X"A7",X"18",X"19",X"CB",X"E7",X"16",
		X"02",X"16",X"CB",X"E6",X"18",X"19",X"CB",X"E9",
		X"03",X"1A",X"17",X"1B",X"00",X"00",X"02",X"16",
		X"00",X"03",X"CA",X"17",X"03",X"00",X"19",X"D0",
		X"19",X"C4",X"C5",X"01",X"FF",X"00",X"19",X"CA",
		X"03",X"00",X"19",X"D0",X"19",X"C3",X"C5",X"FF",
		X"CB",X"F5",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"24",X"25",X"00",X"11",X"00",X"19",X"19",X"18",
		X"06",X"18",X"24",X"01",X"24",X"00",X"03",X"CB",
		X"EF",X"26",X"00",X"00",X"27",X"00",X"00",X"28",
		X"00",X"00",X"29",X"00",X"00",X"2A",X"00",X"00",
		X"2B",X"18",X"19",X"26",X"00",X"27",X"00",X"28",
		X"00",X"29",X"00",X"2A",X"00",X"2B",X"00",X"24",
		X"06",X"24",X"19",X"01",X"19",X"16",X"02",X"16",
		X"03",X"CB",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"24",X"25",X"00",X"51",X"00",X"19",X"19",X"18",
		X"06",X"18",X"24",X"01",X"24",X"00",X"03",X"CB",
		X"EF",X"2B",X"00",X"00",X"2A",X"00",X"00",X"29",
		X"00",X"00",X"28",X"00",X"00",X"27",X"00",X"00",
		X"18",X"19",X"00",X"27",X"00",X"28",X"00",X"29",
		X"00",X"2A",X"00",X"2B",X"00",X"24",X"06",X"24",
		X"19",X"01",X"19",X"16",X"02",X"16",X"03",X"CB",
		X"E1",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"24",X"25",X"00",X"93",X"00",X"FF",X"01",X"19",
		X"19",X"18",X"06",X"18",X"24",X"01",X"24",X"00",
		X"03",X"CB",X"EE",X"26",X"00",X"00",X"27",X"00",
		X"00",X"28",X"00",X"00",X"29",X"00",X"00",X"2A",
		X"00",X"00",X"2B",X"18",X"19",X"26",X"00",X"27",
		X"00",X"28",X"00",X"29",X"00",X"2A",X"00",X"2B",
		X"00",X"24",X"06",X"24",X"19",X"01",X"19",X"16",
		X"02",X"16",X"03",X"CB",X"E0",X"00",X"00",X"00",
		X"24",X"25",X"00",X"D3",X"00",X"FF",X"01",X"19",
		X"19",X"18",X"06",X"18",X"24",X"01",X"24",X"00",
		X"03",X"CB",X"EE",X"2B",X"00",X"00",X"2A",X"00",
		X"00",X"29",X"00",X"00",X"28",X"00",X"00",X"27",
		X"00",X"00",X"18",X"19",X"00",X"27",X"00",X"28",
		X"00",X"29",X"00",X"2A",X"00",X"2B",X"00",X"24",
		X"06",X"24",X"19",X"01",X"19",X"16",X"02",X"16",
		X"03",X"CB",X"E1",X"18",X"18",X"01",X"F8",X"19",
		X"00",X"27",X"05",X"05",X"25",X"27",X"03",X"CB",
		X"EF",X"F8",X"28",X"24",X"25",X"00",X"1D",X"28",
		X"00",X"00",X"00",X"0F",X"17",X"17",X"01",X"00",
		X"1D",X"1D",X"1D",X"28",X"00",X"00",X"00",X"0F",
		X"23",X"23",X"01",X"00",X"1D",X"1D",X"1D",X"28",
		X"00",X"00",X"00",X"0F",X"2F",X"2F",X"01",X"00",
		X"1D",X"1D",X"1D",X"28",X"00",X"00",X"00",X"0F",
		X"3B",X"3B",X"01",X"00",X"1D",X"1D",X"1D",X"28",
		X"00",X"00",X"00",X"0F",X"47",X"47",X"01",X"00",
		X"1D",X"1D",X"1D",X"28",X"00",X"00",X"00",X"0F",
		X"53",X"53",X"01",X"00",X"1D",X"1D",X"1D",X"28",
		X"00",X"00",X"00",X"0F",X"5F",X"5F",X"01",X"00",
		X"1D",X"1D",X"1D",X"28",X"00",X"00",X"00",X"0F",
		X"6B",X"6B",X"01",X"00",X"1D",X"1D",X"24",X"27",
		X"00",X"24",X"01",X"24",X"26",X"7C",X"16",X"02",
		X"16",X"03",X"00",X"BD",X"03",X"00",X"BE",X"05",
		X"F5",X"FF",X"15",X"25",X"FC",X"15",X"9A",X"27",
		X"01",X"7F",X"80",X"19",X"27",X"FE",X"27",X"00",
		X"01",X"27",X"27",X"EE",X"1D",X"00",X"FE",X"05",
		X"00",X"FF",X"0E",X"F2",X"F6",X"25",X"27",X"FE",
		X"27",X"00",X"01",X"27",X"27",X"E7",X"1D",X"00",
		X"FE",X"05",X"00",X"FF",X"25",X"00",X"80",X"1D",
		X"27",X"01",X"00",X"00",X"00",X"28",X"29",X"27",
		X"FE",X"1D",X"00",X"27",X"0E",X"F0",X"20",X"25",
		X"00",X"80",X"1D",X"B2",X"00",X"00",X"24",X"1A",
		X"25",X"1B",X"0E",X"20",X"F6",X"00",X"25",X"00",
		X"00",X"1A",X"00",X"1B",X"0E",X"20",X"F5",X"1C",
		X"00",X"01",X"1C",X"00",X"18",X"28",X"29",X"0E",
		X"F4",X"20",X"0E",X"1C",X"01",X"1C",X"18",X"00",
		X"20",X"F6",X"02",X"05",X"00",X"19",X"03",X"FB",
		X"CB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",
		X"06",X"E0",X"42",X"58",X"5D",X"5D",X"5D",X"58",
		X"58",X"42",X"52",X"58",X"78",X"78",X"78",X"58",
		X"CF",X"AB",X"42",X"58",X"5B",X"5B",X"5B",X"58",
		X"58",X"7B",X"58",X"58",X"7A",X"7A",X"7A",X"58",
		X"15",X"3A",X"15",X"1A",X"1B",X"00",X"26",X"1A",
		X"01",X"1A",X"2D",X"2E",X"00",X"01",X"1B",X"1B",
		X"26",X"1F",X"00",X"34",X"00",X"26",X"45",X"1B",
		X"F2",X"F3",X"13",X"3B",X"01",X"0D",X"05",X"01",
		X"1E",X"00",X"00",X"00",X"1B",X"25",X"1A",X"24",
		X"01",X"1A",X"4D",X"4E",X"00",X"01",X"1B",X"1B",
		X"F2",X"EE",X"18",X"24",X"00",X"25",X"F2",X"F2",
		X"00",X"F2",X"F4",X"5F",X"2A",X"5F",X"00",X"24",
		X"00",X"25",X"01",X"1A",X"1A",X"68",X"69",X"00",
		X"01",X"1B",X"1B",X"F2",X"EE",X"70",X"71",X"00",
		X"FF",X"1B",X"1B",X"1A",X"01",X"1A",X"20",X"ED",
		X"7D",X"00",X"7D",X"2A",X"2B",X"24",X"F3",X"15",
		X"6D",X"1A",X"26",X"BE",X"87",X"88",X"24",X"2B",
		X"00",X"24",X"8E",X"00",X"90",X"00",X"00",X"00",
		X"80",X"00",X"25",X"1A",X"01",X"1A",X"99",X"9A",
		X"00",X"01",X"1B",X"1B",X"00",X"25",X"25",X"1A",
		X"01",X"1A",X"A5",X"A6",X"00",X"01",X"1B",X"1B",
		X"24",X"F2",X"E0",X"00",X"00",X"F8",X"15",X"00",
		X"6D",X"1A",X"01",X"1A",X"B7",X"B8",X"00",X"01",
		X"1B",X"1B",X"00",X"00",X"24",X"00",X"25",X"2B",
		X"24",X"24",X"C6",X"2B",X"C8",X"2B",X"2B",X"00",
		X"80",X"00",X"25",X"25",X"24",X"F2",X"E5",X"24",
		X"D3",X"D4",X"00",X"FF",X"25",X"1A",X"01",X"1A",
		X"DB",X"DC",X"00",X"01",X"1B",X"1B",X"F2",X"EE",
		X"2A",X"1D",X"01",X"00",X"25",X"1D",X"00",X"24",
		X"1A",X"01",X"1A",X"EE",X"EF",X"00",X"01",X"1B",
		X"1B",X"ED",X"15",X"F8",X"15",X"0F",X"26",X"FF",
		X"13",X"F9",X"01",X"10",X"05",X"01",X"1E",X"00",
		X"FD",X"89",X"FD",X"FD",X"FD",X"89",X"F1",X"FD",
		X"F3",X"89",X"F1",X"FD",X"FD",X"89",X"F1",X"FD",
		X"3F",X"89",X"FD",X"FD",X"FD",X"89",X"F1",X"FD",
		X"36",X"89",X"FD",X"FD",X"FD",X"89",X"F1",X"FD",
		X"9A",X"85",X"FD",X"FD",X"F5",X"85",X"F7",X"FD",
		X"F9",X"85",X"F7",X"FD",X"F5",X"85",X"F7",X"FD",
		X"42",X"85",X"FD",X"FD",X"FD",X"85",X"F7",X"FD",
		X"38",X"85",X"FD",X"FD",X"FD",X"85",X"F7",X"FD",
		X"D3",X"8C",X"FD",X"FD",X"FD",X"8C",X"D7",X"FD",
		X"D9",X"8C",X"D7",X"FD",X"96",X"8C",X"D7",X"FD",
		X"45",X"8C",X"FD",X"FD",X"FD",X"8C",X"D7",X"FD",
		X"DB",X"8C",X"FD",X"FD",X"FD",X"8C",X"D7",X"FD",
		X"DD",X"01",X"FD",X"FD",X"FD",X"01",X"D5",X"FD",
		X"DF",X"01",X"D5",X"FD",X"98",X"01",X"D5",X"FD",
		X"49",X"01",X"FD",X"FD",X"FD",X"01",X"D5",X"FD",
		X"E1",X"01",X"FD",X"FD",X"FD",X"01",X"D5",X"FD",
		X"FD",X"C1",X"FD",X"FD",X"C7",X"C1",X"C3",X"FD",
		X"7F",X"FD",X"CD",X"FD",X"C7",X"C1",X"C3",X"FD",
		X"4D",X"C1",X"FD",X"FD",X"C7",X"C1",X"C5",X"FD",
		X"CF",X"C1",X"E3",X"FD",X"FD",X"C1",X"FD",X"FD",
		X"BF",X"B9",X"BB",X"FD",X"BF",X"B9",X"BB",X"FD",
		X"CB",X"B9",X"C9",X"FD",X"BF",X"B9",X"BB",X"FD",
		X"51",X"B9",X"FD",X"FD",X"BF",X"B9",X"BD",X"FD",
		X"D1",X"B9",X"E5",X"FD",X"BF",X"B9",X"BB",X"FD",
		X"E7",X"E9",X"FD",X"FD",X"E7",X"E9",X"EB",X"FD",
		X"7B",X"E9",X"77",X"FD",X"E7",X"E9",X"EB",X"FD",
		X"55",X"E9",X"FD",X"FD",X"FD",X"E9",X"EB",X"FD",
		X"ED",X"E9",X"FD",X"FD",X"FD",X"E9",X"EB",X"FD",
		X"EF",X"29",X"FD",X"FD",X"EF",X"29",X"B7",X"FD",
		X"6C",X"29",X"83",X"FD",X"EF",X"29",X"B7",X"FD",
		X"58",X"29",X"FD",X"FD",X"FD",X"29",X"B7",X"FD",
		X"FB",X"29",X"FD",X"FD",X"FD",X"29",X"B7",X"00",
		X"0E",X"25",X"27",X"18",X"20",X"00",X"28",X"29",
		X"18",X"18",X"00",X"28",X"18",X"80",X"1D",X"28",
		X"18",X"15",X"00",X"17",X"00",X"00",X"00",X"80",
		X"27",X"7E",X"00",X"1D",X"27",X"0E",X"20",X"ED",
		X"18",X"28",X"29",X"27",X"7F",X"27",X"0E",X"F4",
		X"20",X"25",X"00",X"FF",X"19",X"19",X"24",X"00",
		X"25",X"69",X"26",X"0E",X"F2",X"F5",X"27",X"3B",
		X"FE",X"27",X"01",X"27",X"00",X"20",X"F8",X"29",
		X"75",X"5B",X"29",X"75",X"5B",X"27",X"80",X"5B",
		X"3D",X"27",X"80",X"5B",X"3D",X"27",X"01",X"5B",
		X"3D",X"27",X"01",X"5B",X"3D",X"28",X"75",X"5B",
		X"28",X"75",X"5B",X"24",X"1A",X"1A",X"62",X"24",
		X"64",X"24",X"24",X"00",X"80",X"00",X"25",X"1B",
		X"1B",X"00",X"20",X"F2",X"00",X"2A",X"01",X"2A",
		X"28",X"29",X"F7",X"20",X"00",X"20",X"F9",X"2A",
		X"01",X"70",X"2A",X"2B",X"01",X"70",X"2B",X"2B",
		X"01",X"70",X"2B",X"FA",X"20",X"25",X"18",X"90",
		X"00",X"25",X"18",X"90",X"00",X"25",X"18",X"00",
		X"18",X"28",X"29",X"0E",X"F6",X"20",X"0D",X"C5",
		X"0D",X"CD",X"1C",X"02",X"1C",X"00",X"1B",X"25",
		X"1A",X"24",X"01",X"1A",X"00",X"A8",X"A9",X"00",
		X"01",X"1B",X"1B",X"00",X"24",X"25",X"00",X"1A",
		X"1A",X"1B",X"00",X"1B",X"0E",X"ED",X"20",X"11",
		X"0E",X"11",X"18",X"11",X"22",X"11",X"2A",X"11",
		X"26",X"11",X"34",X"11",X"3A",X"11",X"40",X"11",
		X"48",X"11",X"4D",X"11",X"62",X"11",X"65",X"11",
		X"68",X"11",X"76",X"11",X"E4",X"0D",X"83",X"0D",
		X"9D",X"0D",X"E2",X"11",X"6B",X"11",X"8F",X"0D",
		X"D7",X"11",X"6E",X"11",X"5E",X"11",X"54",X"11",
		X"BD",X"11",X"BE",X"11",X"05",X"11",X"71",X"11",
		X"BB",X"0D",X"BF",X"11",X"A2",X"11",X"7D",X"0D",
		X"AC",X"11",X"D4",X"11",X"74",X"0D",X"EA",X"06",
		X"15",X"24",X"0F",X"26",X"FF",X"25",X"00",X"01",
		X"00",X"28",X"29",X"0E",X"F5",X"20",X"25",X"00",
		X"01",X"00",X"28",X"29",X"0E",X"F5",X"20",X"00",
		X"00",X"25",X"00",X"18",X"28",X"29",X"00",X"0E",
		X"20",X"F5",X"25",X"00",X"1C",X"2A",X"25",X"00",
		X"1C",X"2B",X"24",X"2A",X"2B",X"00",X"2A",X"28",
		X"29",X"0E",X"20",X"F5",X"25",X"18",X"00",X"0E",
		X"20",X"F7",X"25",X"2A",X"00",X"0E",X"20",X"F7",
		X"24",X"2A",X"2B",X"2A",X"00",X"0E",X"20",X"F6",
		X"25",X"2B",X"00",X"0E",X"20",X"F7",X"18",X"2A",
		X"28",X"29",X"0E",X"20",X"F6",X"1C",X"01",X"2A",
		X"28",X"29",X"00",X"0E",X"20",X"F5",X"2A",X"01",
		X"58",X"1C",X"18",X"50",X"2B",X"2A",X"50",X"18",
		X"2B",X"50",X"18",X"27",X"79",X"FB",X"27",X"79",
		X"04",X"27",X"79",X"F7",X"27",X"79",X"08",X"27",
		X"7F",X"27",X"0E",X"F6",X"20",X"00",X"24",X"25",
		X"00",X"29",X"18",X"28",X"27",X"7F",X"27",X"00",
		X"00",X"80",X"27",X"27",X"0E",X"20",X"F1",X"1C",
		X"00",X"02",X"1C",X"00",X"00",X"00",X"01",X"1A",
		X"9B",X"9C",X"00",X"01",X"00",X"1B",X"00",X"0E",
		X"20",X"F1",X"1C",X"01",X"1C",X"27",X"BD",X"AA",
		X"AA",X"C0",X"00",X"28",X"AF",X"B0",X"00",X"02",
		X"00",X"00",X"29",X"80",X"00",X"20",X"00",X"00",
		X"0E",X"20",X"EE",X"C0",X"2A",X"C0",X"2B",X"18",
		X"25",X"C7",X"00",X"28",X"29",X"CB",X"00",X"28",
		X"29",X"00",X"00",X"80",X"80",X"27",X"FE",X"00",
		X"27",X"0E",X"20",X"F1",X"1C",X"00",X"01",X"1C",
		X"00",X"29",X"02",X"02",X"28",X"00",X"7F",X"40",
		X"27",X"0E",X"20",X"F2",X"1C",X"00",X"03",X"1C",
		X"00",X"29",X"02",X"02",X"28",X"00",X"00",X"00",
		X"7F",X"40",X"27",X"00",X"00",X"1A",X"00",X"1B",
		X"00",X"0E",X"20",X"EE",X"00",X"00",X"00",X"00",
		X"F6",X"F7",X"09",X"16",X"55",X"1E",X"05",X"FF",
		X"1F",X"30",X"17",X"31",X"18",X"32",X"19",X"33",
		X"F6",X"02",X"16",X"F7",X"17",X"05",X"19",X"00",
		X"18",X"02",X"05",X"55",X"1E",X"05",X"FF",X"16",
		X"00",X"05",X"30",X"16",X"31",X"17",X"32",X"18",
		X"33",X"19",X"00",X"03",X"0C",X"15",X"0F",X"01",
		X"0F",X"42",X"0F",X"01",X"10",X"39",X"FE",X"00",
		X"3C",X"0F",X"11",X"11",X"0F",X"11",X"11",X"0F",
		X"B3",X"10",X"FF",X"10",X"0F",X"11",X"0F",X"00",
		X"00",X"3E",X"00",X"17",X"1C",X"37",X"1D",X"FE",
		X"16",X"75",X"CF",X"23",X"00",X"5E",X"27",X"CF",
		X"00",X"5E",X"26",X"CF",X"00",X"5E",X"28",X"CF",
		X"00",X"F0",X"26",X"93",X"26",X"1A",X"28",X"E6",
		X"01",X"35",X"72",X"E8",X"00",X"CF",X"18",X"00",
		X"35",X"72",X"E0",X"00",X"63",X"FF",X"22",X"00",
		X"00",X"1A",X"24",X"8C",X"FB",X"35",X"72",X"09",
		X"00",X"5E",X"24",X"93",X"25",X"21",X"24",X"7F",
		X"00",X"93",X"24",X"FF",X"03",X"CB",X"D4",X"00",
		X"1D",X"29",X"26",X"96",X"97",X"24",X"25",X"00",
		X"26",X"00",X"26",X"1D",X"29",X"01",X"26",X"A2",
		X"A3",X"24",X"25",X"00",X"26",X"00",X"26",X"1D",
		X"06",X"90",X"08",X"03",X"CB",X"C2",X"18",X"00",
		X"00",X"18",X"00",X"20",X"B7",X"18",X"B9",X"18",
		X"7F",X"00",X"18",X"20",X"BF",X"C0",X"00",X"3F",
		X"00",X"18",X"00",X"01",X"18",X"40",X"C9",X"CA",
		X"FE",X"00",X"16",X"16",X"03",X"CB",X"E7",X"18",
		X"00",X"1D",X"19",X"00",X"18",X"00",X"00",X"00",
		X"18",X"18",X"19",X"1D",X"00",X"19",X"04",X"19",
		X"E3",X"E4",X"FE",X"00",X"16",X"16",X"03",X"00",
		X"EA",X"30",X"25",X"1A",X"24",X"00",X"26",X"24",
		X"01",X"24",X"00",X"25",X"00",X"25",X"01",X"25",
		X"26",X"EE",X"01",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"BA",X"BE",X"FF",X"FF",X"FE",
		X"EB",X"FF",X"FE",X"FB",X"FB",X"BF",X"FF",X"FA",
		X"AF",X"FF",X"FF",X"AE",X"EF",X"BA",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"EB",X"BF",X"EE",X"EF",X"FE",
		X"AE",X"FF",X"FE",X"EE",X"AF",X"FF",X"FF",X"FF",
		X"FF",X"AF",X"FF",X"FF",X"EF",X"FF",X"BF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"BB",X"BE",X"EB",X"FF",
		X"FA",X"FF",X"BF",X"6F",X"EA",X"BB",X"5A",X"A9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"AF",X"FE",X"FF",X"FF",X"FF",
		X"BF",X"FF",X"FF",X"BB",X"FA",X"FF",X"FF",X"BF",
		X"FA",X"FF",X"FF",X"EB",X"BB",X"BE",X"FF",X"BF",
		X"FF",X"FF",X"FF",X"BE",X"EB",X"FB",X"AF",X"9A",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",
		X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"BB",X"BA",
		X"AA",X"BA",X"FA",X"FF",X"FF",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FE",X"FF",X"FB",X"FF",X"EF",
		X"AB",X"AA",X"FB",X"EF",X"BB",X"BE",X"EB",X"FF",
		X"FF",X"FF",X"BF",X"AE",X"EB",X"FF",X"BF",X"FF",
		X"FF",X"BF",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"EF",X"6A",X"49",X"96",X"10",
		X"08",X"41",X"15",X"55",X"96",X"AA",X"AA",X"AB",
		X"6A",X"5A",X"56",X"65",X"A9",X"EA",X"AA",X"AA",
		X"FF",X"FF",X"AE",X"EB",X"BF",X"BE",X"BF",X"FF",
		X"FF",X"FF",X"FB",X"AA",X"EF",X"AF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"BE",X"9A",X"92",X"24",X"48",X"92",X"10",X"09",
		X"92",X"20",X"08",X"41",X"10",X"04",X"41",X"10",
		X"04",X"41",X"10",X"04",X"42",X"10",X"54",X"AA",
		X"E9",X"FF",X"EB",X"EF",X"FF",X"EB",X"FF",X"FF",
		X"FF",X"FE",X"FF",X"FF",X"FF",X"BF",X"EB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E6",
		X"28",X"4A",X"92",X"24",X"49",X"92",X"20",X"49",
		X"82",X"24",X"08",X"42",X"10",X"04",X"42",X"10",
		X"08",X"81",X"20",X"04",X"81",X"10",X"09",X"91",
		X"50",X"F9",X"EF",X"FF",X"FF",X"FF",X"FF",X"BF",
		X"FF",X"FF",X"EE",X"EF",X"BF",X"BF",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DF",X"E3",
		X"28",X"8F",X"E3",X"28",X"4A",X"92",X"28",X"4D",
		X"92",X"20",X"49",X"82",X"24",X"48",X"82",X"10",
		X"09",X"92",X"24",X"08",X"91",X"24",X"48",X"82",
		X"24",X"55",X"A6",X"BF",X"FF",X"FF",X"FA",X"EF",
		X"BF",X"FF",X"FF",X"AB",X"FF",X"EE",X"EE",X"EA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"9F",X"F2",
		X"3D",X"DB",X"A3",X"38",X"89",X"93",X"24",X"85",
		X"92",X"24",X"49",X"92",X"24",X"09",X"92",X"24",
		X"48",X"92",X"20",X"09",X"92",X"20",X"09",X"41",
		X"20",X"04",X"41",X"E5",X"FF",X"AB",X"FF",X"BF",
		X"9B",X"FA",X"AE",X"EF",X"AA",X"AE",X"EE",X"EA",
		X"FF",X"FF",X"FF",X"FF",X"AF",X"FF",X"FF",X"F7",
		X"69",X"CF",X"F7",X"69",X"56",X"51",X"15",X"11",
		X"10",X"14",X"85",X"92",X"24",X"09",X"92",X"20",
		X"48",X"92",X"24",X"8D",X"92",X"24",X"49",X"42",
		X"10",X"04",X"52",X"10",X"A4",X"FB",X"BB",X"AF",
		X"AB",X"A6",X"59",X"AA",X"BB",X"BA",X"EF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"FE",X"AB",
		X"44",X"DA",X"F7",X"29",X"10",X"50",X"44",X"55",
		X"41",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"04",X"44",X"50",X"24",X"49",X"92",X"24",X"49",
		X"92",X"24",X"89",X"E2",X"34",X"4A",X"92",X"24",
		X"09",X"91",X"24",X"09",X"52",X"BB",X"BF",X"EB",
		X"BA",X"6E",X"97",X"A5",X"59",X"EA",X"FF",X"FF",
		X"EF",X"BF",X"FA",X"EF",X"FE",X"FF",X"AB",X"80",
		X"10",X"A5",X"7D",X"4A",X"11",X"01",X"55",X"11",
		X"15",X"11",X"40",X"14",X"48",X"91",X"20",X"49",
		X"92",X"34",X"09",X"92",X"24",X"08",X"92",X"24",
		X"89",X"93",X"24",X"48",X"96",X"BE",X"FF",X"BF",
		X"BB",X"BF",X"EB",X"A6",X"A9",X"FF",X"FF",X"FF",
		X"FF",X"FA",X"BF",X"FB",X"EB",X"FF",X"A7",X"80",
		X"40",X"54",X"AA",X"4A",X"45",X"80",X"40",X"40",
		X"80",X"00",X"51",X"24",X"49",X"96",X"24",X"49",
		X"D2",X"24",X"49",X"82",X"50",X"89",X"E2",X"28",
		X"49",X"92",X"28",X"49",X"42",X"41",X"F9",X"FB",
		X"FA",X"FB",X"EB",X"FF",X"AE",X"AA",X"FA",X"FF",
		X"FF",X"FF",X"FB",X"FF",X"FF",X"BF",X"57",X"40",
		X"40",X"01",X"41",X"E5",X"AA",X"15",X"51",X"50",
		X"40",X"10",X"00",X"01",X"01",X"51",X"24",X"49",
		X"51",X"24",X"48",X"A2",X"25",X"49",X"92",X"38",
		X"8A",X"A3",X"24",X"49",X"92",X"24",X"49",X"01",
		X"01",X"44",X"55",X"A5",X"BF",X"EB",X"BF",X"AE",
		X"56",X"66",X"F4",X"FF",X"BF",X"BF",X"FF",X"BF",
		X"FE",X"FF",X"15",X"15",X"40",X"95",X"EA",X"57",
		X"40",X"00",X"01",X"02",X"01",X"08",X"04",X"09",
		X"52",X"24",X"09",X"52",X"24",X"49",X"92",X"38",
		X"8A",X"E3",X"28",X"8E",X"93",X"28",X"49",X"92",
		X"10",X"05",X"01",X"01",X"44",X"A6",X"65",X"AA",
		X"EA",X"BA",X"69",X"EA",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"9F",X"41",X"54",X"95",X"FE",
		X"BB",X"5F",X"00",X"03",X"04",X"0C",X"10",X"45",
		X"92",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"24",X"49",X"92",X"24",X"89",X"92",X"24",X"49",
		X"E2",X"28",X"59",X"E2",X"28",X"49",X"11",X"40",
		X"40",X"91",X"24",X"4A",X"92",X"10",X"54",X"EA",
		X"B6",X"AE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"BF",X"4A",X"55",X"95",X"DA",X"A7",X"7F",
		X"05",X"0C",X"05",X"51",X"41",X"14",X"45",X"92",
		X"24",X"8A",X"E2",X"28",X"4E",X"A2",X"24",X"49",
		X"A2",X"24",X"89",X"A2",X"64",X"8A",X"42",X"40",
		X"00",X"61",X"28",X"8E",X"92",X"14",X"54",X"A6",
		X"BB",X"AE",X"FE",X"FF",X"FF",X"FF",X"FF",X"AF",
		X"FE",X"FF",X"5F",X"52",X"59",X"9F",X"AA",X"A9",
		X"AA",X"56",X"15",X"10",X"50",X"40",X"40",X"51",
		X"24",X"49",X"A2",X"38",X"89",X"E2",X"28",X"8A",
		X"92",X"64",X"8F",X"A3",X"28",X"9E",X"56",X"28",
		X"4A",X"52",X"40",X"00",X"A1",X"39",X"8A",X"92",
		X"24",X"45",X"99",X"BA",X"FD",X"FF",X"FF",X"FF",
		X"FF",X"BF",X"AF",X"FE",X"FF",X"9B",X"A6",X"A9",
		X"A6",X"BE",X"BA",X"EB",X"AB",X"6A",X"55",X"A1",
		X"24",X"49",X"A6",X"28",X"8A",X"92",X"68",X"8E",
		X"A3",X"78",X"9B",X"F3",X"39",X"4A",X"56",X"14",
		X"89",X"92",X"24",X"04",X"04",X"14",X"8A",X"A6",
		X"28",X"4A",X"96",X"94",X"FE",X"FF",X"BF",X"FE",
		X"FF",X"FF",X"BF",X"FB",X"FB",X"9F",X"96",X"64",
		X"DA",X"EB",X"FE",X"EB",X"AF",X"FE",X"EF",X"A7",
		X"28",X"8A",X"A2",X"24",X"8A",X"E3",X"39",X"CE",
		X"F2",X"38",X"8E",X"FA",X"7A",X"5A",X"52",X"28",
		X"49",X"91",X"28",X"49",X"42",X"14",X"89",X"A2",
		X"28",X"45",X"66",X"24",X"AA",X"57",X"95",X"59",
		X"99",X"FF",X"FF",X"FF",X"2A",X"49",X"91",X"28",
		X"99",X"B3",X"79",X"EA",X"FB",X"AE",X"DE",X"A3",
		X"78",X"8A",X"E2",X"28",X"CE",X"A3",X"3C",X"9A",
		X"F3",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"29",X"9E",X"F6",X"28",X"8A",X"92",X"28",X"8E",
		X"92",X"28",X"8A",X"92",X"24",X"8A",X"B7",X"28",
		X"89",X"92",X"29",X"99",X"96",X"A2",X"59",X"9A",
		X"FF",X"FF",X"A7",X"14",X"44",X"92",X"28",X"8A",
		X"A2",X"28",X"9A",X"FA",X"7D",X"9F",X"A3",X"7E",
		X"8E",X"A2",X"68",X"DA",X"A3",X"79",X"8F",X"A3",
		X"38",X"CA",X"A3",X"38",X"8A",X"E6",X"28",X"8E",
		X"E2",X"38",X"8E",X"E2",X"28",X"8A",X"F6",X"28",
		X"8A",X"92",X"24",X"4A",X"DA",X"A6",X"BE",X"FF",
		X"FF",X"9F",X"42",X"24",X"49",X"91",X"28",X"DE",
		X"A7",X"68",X"9A",X"F6",X"AD",X"EF",X"FB",X"BE",
		X"9F",X"E2",X"6D",X"DF",X"A7",X"7D",X"DF",X"A3",
		X"7D",X"9F",X"F7",X"28",X"9E",X"F3",X"7D",X"DE",
		X"B3",X"39",X"8A",X"A3",X"24",X"4A",X"A2",X"38",
		X"9A",X"A2",X"64",X"AA",X"EB",X"BA",X"FA",X"FF",
		X"FF",X"4F",X"A1",X"29",X"89",X"A2",X"39",X"9A",
		X"EA",X"69",X"AA",X"F7",X"B9",X"EF",X"AB",X"BE",
		X"9F",X"F6",X"7D",X"DE",X"F7",X"7D",X"EF",X"F7",
		X"7D",X"DF",X"F7",X"7D",X"DF",X"B7",X"39",X"8B",
		X"E3",X"28",X"8E",X"E2",X"28",X"8A",X"A3",X"6D",
		X"8A",X"A2",X"68",X"A9",X"AA",X"AA",X"AA",X"EF",
		X"7E",X"45",X"A5",X"28",X"9A",X"F6",X"69",X"8B",
		X"F6",X"AA",X"EF",X"FB",X"BE",X"DE",X"FB",X"BD",
		X"EF",X"E7",X"6E",X"EF",X"F7",X"BE",X"9F",X"F7",
		X"79",X"DA",X"FB",X"79",X"8F",X"E3",X"28",X"8E",
		X"E2",X"28",X"8A",X"A3",X"28",X"8A",X"E2",X"78",
		X"5F",X"E6",X"28",X"69",X"9A",X"62",X"15",X"A9",
		X"29",X"99",X"E6",X"28",X"4A",X"A2",X"68",X"DE",
		X"E7",X"BD",X"EE",X"FB",X"69",X"DF",X"E7",X"AD",
		X"EE",X"F7",X"BD",X"DF",X"EB",X"6D",X"EF",X"F7",
		X"7D",X"DF",X"A3",X"3D",X"8A",X"E2",X"2C",X"8E",
		X"A2",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"3C",X"8A",X"A3",X"38",X"8E",X"A3",X"68",X"9F",
		X"1A",X"69",X"A5",X"9A",X"BA",X"BE",X"EB",X"66",
		X"DA",X"A3",X"28",X"8A",X"A2",X"68",X"DE",X"A7",
		X"6C",X"EE",X"F7",X"BD",X"9F",X"FB",X"BE",X"EF",
		X"F6",X"7A",X"9B",X"FB",X"7D",X"DE",X"F7",X"6D",
		X"9E",X"E3",X"28",X"DE",X"E2",X"68",X"8F",X"F2",
		X"28",X"8E",X"A2",X"29",X"DF",X"E2",X"68",X"EF",
		X"6B",X"86",X"A6",X"96",X"A6",X"FE",X"EE",X"39",
		X"8A",X"92",X"68",X"8E",X"E6",X"68",X"DA",X"F7",
		X"78",X"DA",X"FB",X"79",X"EF",X"F6",X"BE",X"EF",
		X"FB",X"7D",X"DF",X"F6",X"79",X"DF",X"E6",X"7D",
		X"DF",X"B7",X"7C",X"8F",X"F3",X"38",X"8A",X"B3",
		X"38",X"8A",X"E2",X"68",X"CF",X"E7",X"BD",X"9B",
		X"6B",X"85",X"A5",X"99",X"55",X"A4",X"FB",X"64",
		X"56",X"A2",X"69",X"DE",X"B3",X"78",X"9A",X"B7",
		X"7D",X"DF",X"F7",X"BD",X"EF",X"EB",X"FE",X"EF",
		X"E7",X"6E",X"EE",X"F7",X"69",X"DF",X"F7",X"3D",
		X"DE",X"F7",X"79",X"DB",X"B3",X"38",X"8B",X"E2",
		X"28",X"8F",X"E2",X"78",X"8B",X"B3",X"7D",X"DE",
		X"6B",X"86",X"A6",X"DA",X"A6",X"FA",X"FE",X"65",
		X"A1",X"F9",X"7E",X"DA",X"A3",X"68",X"9F",X"E6",
		X"B9",X"EE",X"B7",X"7A",X"EF",X"FB",X"FF",X"DB",
		X"BB",X"39",X"DF",X"A7",X"3C",X"DA",X"E3",X"7D",
		X"9B",X"B7",X"3D",X"DF",X"E3",X"2D",X"8E",X"F7",
		X"78",X"8F",X"E2",X"69",X"8F",X"A2",X"7C",X"DA",
		X"AB",X"86",X"A6",X"E9",X"A6",X"6E",X"AA",X"9A",
		X"A1",X"A6",X"68",X"9F",X"A2",X"A8",X"9E",X"F6",
		X"78",X"9F",X"F7",X"7E",X"9F",X"FA",X"7E",X"EE",
		X"A6",X"7D",X"DA",X"A3",X"7D",X"8B",X"B7",X"3D",
		X"DF",X"F3",X"3D",X"DA",X"B3",X"3C",X"DE",X"A2",
		X"7C",X"CA",X"F3",X"7D",X"8F",X"A2",X"68",X"8F",
		X"A7",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"8A",X"A6",X"EE",X"BA",X"59",X"55",X"85",X"A6",
		X"A2",X"68",X"CE",X"E6",X"68",X"AE",X"E6",X"AA",
		X"EF",X"B7",X"79",X"DF",X"FB",X"7E",X"9B",X"F7",
		X"39",X"9F",X"E6",X"6C",X"CE",X"F3",X"3D",X"DE",
		X"A3",X"7D",X"CF",X"F7",X"7D",X"CA",X"E3",X"28",
		X"9F",X"A3",X"79",X"8F",X"E2",X"28",X"DA",X"BB",
		X"96",X"AA",X"DA",X"A6",X"6E",X"06",X"86",X"86",
		X"A3",X"29",X"8A",X"F6",X"68",X"AE",X"FB",X"BE",
		X"FE",X"F7",X"BE",X"9F",X"FA",X"7E",X"DF",X"B7",
		X"78",X"DA",X"F3",X"3C",X"CA",X"A7",X"3C",X"DB",
		X"F7",X"7C",X"9B",X"F3",X"68",X"CF",X"A7",X"7C",
		X"CE",X"E2",X"7D",X"8F",X"A2",X"28",X"8E",X"A7",
		X"8A",X"BA",X"9A",X"BA",X"AD",X"17",X"56",X"8A",
		X"A6",X"39",X"8A",X"A3",X"78",X"9A",X"EA",X"BE",
		X"EB",X"EF",X"BE",X"EF",X"FB",X"7D",X"CA",X"E7",
		X"7C",X"8F",X"E2",X"2D",X"DE",X"E2",X"6C",X"8E",
		X"B3",X"39",X"DF",X"F6",X"7C",X"DF",X"F3",X"6D",
		X"8F",X"F7",X"6C",X"DF",X"A3",X"38",X"8B",X"A6",
		X"9A",X"6A",X"FF",X"FF",X"BF",X"16",X"1A",X"4A",
		X"AA",X"29",X"8B",X"A3",X"28",X"AE",X"E6",X"FA",
		X"FF",X"FB",X"BF",X"EB",X"FB",X"79",X"DF",X"B3",
		X"29",X"DE",X"B3",X"38",X"8B",X"F3",X"39",X"DB",
		X"F3",X"3D",X"DE",X"F7",X"29",X"8F",X"F6",X"78",
		X"DF",X"F2",X"39",X"9F",X"F7",X"3D",X"8A",X"A3",
		X"AA",X"BE",X"EB",X"FA",X"FF",X"1B",X"5A",X"8A",
		X"A6",X"39",X"CA",X"E6",X"65",X"9A",X"A7",X"BA",
		X"FE",X"FE",X"FE",X"FF",X"FB",X"7D",X"CE",X"F6",
		X"78",X"8F",X"F6",X"28",X"CE",X"A7",X"6C",X"CE",
		X"A3",X"3D",X"DB",X"B3",X"7D",X"DF",X"F7",X"3D",
		X"9F",X"F7",X"78",X"DB",X"E7",X"2C",X"8E",X"A3",
		X"A9",X"5D",X"9A",X"EA",X"EE",X"1A",X"29",X"9E",
		X"A6",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"28",X"89",X"A7",X"7E",X"99",X"E6",X"AA",X"EF",
		X"EF",X"FF",X"EF",X"B7",X"79",X"CB",X"E3",X"2D",
		X"CE",X"A3",X"7C",X"CA",X"F7",X"7C",X"CF",X"F6",
		X"78",X"DF",X"E7",X"7C",X"9F",X"F2",X"68",X"EF",
		X"F6",X"AC",X"EF",X"FB",X"7E",X"CE",X"A2",X"BA",
		X"5E",X"96",X"A6",X"BE",X"6A",X"78",X"9A",X"E6",
		X"28",X"4A",X"E6",X"69",X"5A",X"96",X"B9",X"FE",
		X"FF",X"FF",X"AF",X"FB",X"3D",X"9F",X"B7",X"38",
		X"9B",X"B3",X"38",X"8A",X"B7",X"78",X"8B",X"F7",
		X"6C",X"CE",X"F6",X"6D",X"DF",X"E3",X"7D",X"EF",
		X"A7",X"B8",X"EF",X"AF",X"FE",X"9F",X"EA",X"FB",
		X"AE",X"A7",X"EA",X"FE",X"6A",X"7D",X"85",X"A2",
		X"28",X"9A",X"AA",X"69",X"9A",X"96",X"B9",X"AA",
		X"FF",X"BF",X"AA",X"A6",X"7D",X"8B",X"F3",X"68",
		X"CF",X"E3",X"2D",X"DE",X"F7",X"3D",X"DB",X"F7",
		X"69",X"DF",X"F7",X"7D",X"DE",X"B7",X"7C",X"EE",
		X"A3",X"BC",X"EE",X"FF",X"BF",X"BA",X"DB",X"BA",
		X"BA",X"9B",X"FA",X"AF",X"6A",X"68",X"8A",X"A2",
		X"38",X"8A",X"EB",X"6A",X"9A",X"A6",X"A5",X"AA",
		X"FB",X"BF",X"9A",X"F7",X"7C",X"CE",X"F6",X"7C",
		X"9F",X"F6",X"28",X"DF",X"B7",X"7C",X"CE",X"E6",
		X"7C",X"DF",X"E7",X"7C",X"CF",X"F7",X"AD",X"FF",
		X"E7",X"AE",X"FE",X"EA",X"E9",X"AE",X"9B",X"BA",
		X"69",X"EA",X"BB",X"AE",X"AA",X"68",X"9A",X"A3",
		X"39",X"AE",X"A6",X"65",X"5A",X"96",X"A9",X"EE",
		X"FF",X"AB",X"DA",X"E7",X"2D",X"8F",X"F7",X"68",
		X"DF",X"FB",X"7E",X"9F",X"F2",X"39",X"DB",X"F3",
		X"2D",X"CE",X"F6",X"2C",X"DE",X"E6",X"FD",X"FF",
		X"FB",X"BF",X"FE",X"EA",X"FA",X"AE",X"9B",X"B6",
		X"BE",X"DB",X"A5",X"1A",X"69",X"39",X"9E",X"A2",
		X"79",X"AA",X"EA",X"A9",X"99",X"A6",X"A5",X"AE",
		X"EB",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"BE",X"9A",X"F3",X"7D",X"DF",X"F2",X"7D",X"EF",
		X"EA",X"6E",X"CF",X"F7",X"6C",X"CE",X"E2",X"38",
		X"8B",X"F3",X"69",X"EF",X"F7",X"FE",X"FF",X"FF",
		X"EA",X"AA",X"AB",X"FF",X"AE",X"97",X"E6",X"FE",
		X"EB",X"76",X"08",X"55",X"7F",X"9A",X"E2",X"79",
		X"59",X"EA",X"6A",X"5A",X"96",X"A9",X"AE",X"FB",
		X"7F",X"DE",X"B7",X"39",X"9F",X"F7",X"69",X"55",
		X"55",X"95",X"EA",X"A7",X"7D",X"EF",X"FB",X"AE",
		X"AF",X"BB",X"BE",X"EF",X"F7",X"BE",X"FB",X"AB",
		X"AA",X"BF",X"EF",X"FA",X"FF",X"EB",X"F6",X"EF",
		X"97",X"76",X"59",X"85",X"6A",X"9A",X"A7",X"69",
		X"5A",X"E6",X"BA",X"AA",X"EA",X"A9",X"AE",X"FF",
		X"7F",X"9A",X"F7",X"7D",X"DF",X"A7",X"55",X"95",
		X"55",X"15",X"A5",X"FE",X"BF",X"FA",X"AB",X"AA",
		X"AA",X"AA",X"FF",X"EF",X"EB",X"BE",X"AF",X"AB",
		X"FE",X"BE",X"EB",X"BB",X"FD",X"EF",X"FB",X"BF",
		X"EB",X"76",X"69",X"96",X"BA",X"9A",X"A6",X"65",
		X"85",X"96",X"BA",X"9A",X"AB",X"BA",X"9E",X"AB",
		X"7F",X"DE",X"F7",X"6D",X"9F",X"55",X"99",X"AA",
		X"56",X"45",X"55",X"A9",X"9A",X"AA",X"AA",X"55",
		X"AA",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",
		X"B6",X"AE",X"EF",X"FF",X"AE",X"BF",X"FF",X"FF",
		X"EF",X"BA",X"AE",X"EF",X"7F",X"A5",X"96",X"69",
		X"5A",X"A6",X"A9",X"AF",X"E6",X"B9",X"AA",X"FB",
		X"BF",X"9A",X"E7",X"7A",X"5A",X"55",X"56",X"65",
		X"55",X"55",X"55",X"55",X"A5",X"65",X"A9",X"56",
		X"95",X"55",X"AA",X"A5",X"99",X"9A",X"65",X"55",
		X"56",X"65",X"95",X"AB",X"FE",X"FF",X"FF",X"FF",
		X"AB",X"AA",X"6D",X"FB",X"AF",X"96",X"A6",X"66",
		X"5A",X"A6",X"B9",X"AA",X"AB",X"BA",X"EE",X"FF",
		X"BF",X"6A",X"55",X"55",X"51",X"55",X"95",X"A5",
		X"6A",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"A5",X"A6",X"56",X"9A",X"A9",X"A9",X"6A",X"A5",
		X"9A",X"AA",X"6A",X"A5",X"56",X"6A",X"65",X"56",
		X"A5",X"55",X"56",X"66",X"AA",X"FF",X"FF",X"DB",
		X"BA",X"6E",X"DA",X"BF",X"AA",X"AA",X"6A",X"9A",
		X"A6",X"A5",X"AE",X"E6",X"AA",X"AE",X"6A",X"55",
		X"54",X"54",X"56",X"65",X"59",X"56",X"65",X"A9",
		X"6A",X"E5",X"AF",X"FA",X"EA",X"EB",X"BF",X"5A",
		X"69",X"BF",X"AF",X"BB",X"BB",X"AA",X"AA",X"A6",
		X"66",X"5A",X"95",X"55",X"55",X"A6",X"FA",X"D7",
		X"BA",X"5E",X"97",X"BA",X"AA",X"AA",X"AA",X"9A",
		X"A6",X"A9",X"AE",X"AB",X"65",X"55",X"44",X"45",
		X"65",X"55",X"56",X"65",X"A5",X"AA",X"AA",X"FE",
		X"59",X"A5",X"FE",X"FE",X"AF",X"EA",X"BF",X"9A",
		X"EA",X"BF",X"FB",X"FF",X"BA",X"BE",X"EF",X"BF",
		X"AE",X"AA",X"AA",X"65",X"59",X"99",X"55",X"85",
		X"A6",X"AE",X"97",X"B6",X"5A",X"A9",X"BE",X"6E",
		X"E6",X"6A",X"6A",X"55",X"45",X"51",X"55",X"96",
		X"55",X"59",X"AA",X"AA",X"6A",X"AA",X"AA",X"FE",
		X"6A",X"66",X"F9",X"AB",X"AA",X"AA",X"FF",X"FF",
		X"FE",X"BE",X"FE",X"EB",X"AE",X"6E",X"FB",X"FA",
		X"BE",X"EB",X"BB",X"AE",X"6A",X"66",X"65",X"E9",
		X"F5",X"FE",X"97",X"F5",X"5B",X"55",X"AA",X"EF",
		X"AA",X"55",X"54",X"44",X"95",X"65",X"59",X"A5",
		X"A6",X"A6",X"69",X"EF",X"AB",X"AA",X"EA",X"EA",
		X"FA",X"AF",X"AA",X"6A",X"B5",X"FE",X"BF",X"FF",
		X"FB",X"FB",X"EF",X"EB",X"EA",X"FE",X"AF",X"B6",
		X"6E",X"EF",X"B6",X"6E",X"EB",X"AA",X"6A",X"AD",
		X"FF",X"FF",X"EF",X"FF",X"9E",X"56",X"69",X"6A",
		X"45",X"41",X"51",X"59",X"99",X"55",X"6A",X"AA",
		X"AE",X"EA",X"69",X"EE",X"EB",X"9A",X"AA",X"AA",
		X"BA",X"EA",X"AB",X"AA",X"EA",X"FF",X"EA",X"BF",
		X"FB",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"BF",X"EE",X"EA",X"BF",X"FE",X"AB",X"A6",X"A9",
		X"DB",X"B7",X"7E",X"DB",X"F6",X"AF",X"EA",X"BB",
		X"FF",X"FF",X"FE",X"AF",X"56",X"55",X"54",X"10",
		X"95",X"59",X"59",X"56",X"AA",X"FB",X"6A",X"9A",
		X"B6",X"7A",X"EB",X"FF",X"AA",X"A6",X"AA",X"AE",
		X"AA",X"AA",X"9A",X"FA",X"FB",X"FA",X"EF",X"FE",
		X"BE",X"EE",X"FF",X"FF",X"FE",X"EF",X"FE",X"6F",
		X"DB",X"FA",X"FE",X"EB",X"EB",X"FF",X"AB",X"EA",
		X"BA",X"EF",X"AB",X"9A",X"45",X"45",X"50",X"59",
		X"5A",X"65",X"A9",X"FA",X"AF",X"EB",X"BB",X"AB",
		X"EA",X"7D",X"FE",X"FA",X"AA",X"95",X"69",X"A5",
		X"9A",X"5A",X"9A",X"EA",X"AB",X"AA",X"EF",X"FF",
		X"BE",X"FA",X"FF",X"FB",X"FF",X"FF",X"FF",X"BF",
		X"AB",X"E6",X"FF",X"FF",X"FA",X"FF",X"EB",X"EA",
		X"EF",X"EF",X"6A",X"14",X"04",X"55",X"65",X"95",
		X"96",X"AA",X"E7",X"FA",X"EB",X"FF",X"FE",X"9E",
		X"BA",X"B9",X"AF",X"FB",X"6A",X"66",X"55",X"6A",
		X"65",X"55",X"9A",X"AF",X"EA",X"E9",X"BF",X"FB",
		X"EA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"BF",X"EF",X"FF",X"FF",X"EF",X"FB",
		X"FF",X"5B",X"55",X"50",X"54",X"5A",X"69",X"69",
		X"6A",X"AE",X"AB",X"BA",X"FE",X"FF",X"FA",X"9B",
		X"A6",X"79",X"EA",X"AB",X"AA",X"56",X"55",X"99",
		X"95",X"15",X"AA",X"EE",X"A6",X"AA",X"EF",X"AB",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"BF",X"FE",
		X"FF",X"FF",X"EF",X"EF",X"FE",X"BF",X"9B",X"BA",
		X"6E",X"01",X"41",X"50",X"55",X"96",X"55",X"A9",
		X"B9",X"AF",X"EA",X"BE",X"AE",X"BF",X"FA",X"AF",
		X"A6",X"7E",X"DE",X"AB",X"AA",X"9A",X"59",X"95",
		X"55",X"15",X"5A",X"9A",X"AA",X"A9",X"EA",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",X"FF",X"BF",
		X"BF",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"FB",X"FF",X"AF",X"FF",X"FF",X"FB",X"BB",X"5A",
		X"04",X"45",X"A5",X"59",X"56",X"AA",X"E6",X"AD",
		X"EE",X"EB",X"FA",X"AB",X"FB",X"BA",X"AF",X"A6",
		X"69",X"9E",X"F6",X"AA",X"AA",X"55",X"45",X"56",
		X"54",X"6A",X"EA",X"A6",X"A5",X"AB",X"FF",X"BF",
		X"FE",X"FF",X"FF",X"EB",X"EF",X"EF",X"FF",X"FB",
		X"FF",X"EF",X"FF",X"FF",X"FF",X"FF",X"6A",X"10",
		X"54",X"95",X"59",X"59",X"69",X"AA",X"A6",X"B9",
		X"AB",X"BB",X"BA",X"EE",X"AB",X"FE",X"AF",X"A2",
		X"69",X"9A",X"A7",X"BA",X"9A",X"19",X"45",X"55",
		X"A8",X"69",X"9A",X"A6",X"A9",X"69",X"EA",X"A6",
		X"A9",X"EB",X"FB",X"FE",X"FF",X"FF",X"FF",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"45",X"50",
		X"55",X"5A",X"65",X"AA",X"25",X"AA",X"E7",X"A9",
		X"9F",X"BB",X"BA",X"AF",X"FB",X"BA",X"9A",X"92",
		X"69",X"9A",X"A7",X"A9",X"6B",X"65",X"56",X"61",
		X"65",X"69",X"AA",X"A2",X"95",X"6D",X"DB",X"BA",
		X"BE",X"EA",X"BB",X"BE",X"FF",X"FF",X"AF",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"41",X"55",
		X"59",X"96",X"AA",X"EF",X"69",X"AA",X"AA",X"79",
		X"AB",X"AB",X"BD",X"AA",X"FB",X"AB",X"9B",X"56",
		X"39",X"9A",X"E6",X"AA",X"AA",X"55",X"9A",X"96",
		X"66",X"65",X"AA",X"92",X"A9",X"AE",X"FF",X"FF",
		X"EF",X"EF",X"EA",X"FE",X"FB",X"FF",X"FF",X"EF",
		X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"95",X"A5",
		X"56",X"EA",X"BE",X"DA",X"6A",X"9A",X"F7",X"69",
		X"EA",X"B7",X"AA",X"EE",X"EB",X"BE",X"9A",X"96",
		X"68",X"9A",X"A6",X"A9",X"AA",X"55",X"56",X"5A",
		X"A5",X"69",X"9A",X"56",X"9A",X"ED",X"EF",X"AF",
		X"FE",X"EE",X"BA",X"BE",X"FF",X"EA",X"FA",X"FF",
		X"FE",X"FF",X"FB",X"FF",X"FF",X"FF",X"56",X"66",
		X"A9",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"FF",X"FF",X"EB",X"6A",X"AA",X"EA",X"69",X"9A",
		X"AB",X"A9",X"EB",X"EB",X"6E",X"5A",X"A1",X"25",
		X"9A",X"A7",X"65",X"AA",X"25",X"59",X"9A",X"95",
		X"59",X"9A",X"92",X"AA",X"6E",X"EB",X"A6",X"AA",
		X"EB",X"BB",X"AE",X"EE",X"A6",X"BE",X"BF",X"FF",
		X"FE",X"FE",X"FF",X"FF",X"FF",X"A9",X"B5",X"FF",
		X"FF",X"AF",X"EB",X"7B",X"EA",X"A7",X"7A",X"9A",
		X"B7",X"7A",X"AA",X"FE",X"6A",X"5A",X"A5",X"64",
		X"9A",X"A6",X"59",X"EA",X"5A",X"55",X"56",X"66",
		X"65",X"4A",X"56",X"AA",X"BE",X"EB",X"BA",X"AD",
		X"EB",X"FB",X"BE",X"EB",X"FB",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"AE",X"FF",X"00",X"00",X"00",
		X"AA",X"AE",X"AA",X"A5",X"99",X"9B",X"A9",X"A9",
		X"96",X"6A",X"69",X"95",X"96",X"6A",X"AA",X"A6",
		X"5A",X"99",X"9A",X"A9",X"AA",X"AA",X"A5",X"9A",
		X"AA",X"A5",X"5A",X"AA",X"A5",X"AA",X"A6",X"AA",
		X"AA",X"A6",X"56",X"59",X"6A",X"65",X"56",X"66",
		X"55",X"56",X"65",X"69",X"96",X"66",X"A9",X"AA",
		X"6A",X"AE",X"96",X"B9",X"5A",X"96",X"66",X"A9",
		X"96",X"A6",X"99",X"9A",X"A9",X"A5",X"5A",X"A9",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A6",X"6A",X"A9",X"AA",X"A5",
		X"5A",X"5A",X"65",X"55",X"96",X"99",X"AA",X"99",
		X"A9",X"96",X"6A",X"55",X"56",X"69",X"59",X"AA",
		X"BA",X"6A",X"97",X"66",X"59",X"9A",X"69",X"69",
		X"96",X"AA",X"6A",X"69",X"96",X"5A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"A9",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"65",X"55",X"85",X"95",X"6A",X"56",X"55",
		X"59",X"A5",X"A5",X"56",X"AA",X"AA",X"9A",X"66",
		X"5A",X"95",X"95",X"99",X"96",X"A6",X"5A",X"9A",
		X"AA",X"9E",X"9A",X"69",X"59",X"AA",X"A5",X"59",
		X"AA",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"AA",X"AA",X"96",X"AA",X"A5",X"6A",X"A6",X"6A",
		X"AA",X"AA",X"6A",X"59",X"95",X"A5",X"5A",X"56",
		X"55",X"59",X"AA",X"AA",X"9A",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"A9",X"A6",X"AA",X"AA",
		X"AA",X"65",X"69",X"95",X"55",X"A9",X"AA",X"BA",
		X"5A",X"96",X"6A",X"59",X"9A",X"A5",X"AA",X"EA",
		X"AA",X"A9",X"AB",X"BA",X"AA",X"EA",X"AA",X"AA",
		X"EA",X"AA",X"AA",X"AA",X"96",X"6A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AE",X"AA",X"EA",X"AE",X"AA",
		X"BA",X"AA",X"AB",X"AA",X"AA",X"AA",X"AA",X"59",
		X"9A",X"55",X"59",X"96",X"6A",X"69",X"A6",X"A9",
		X"6A",X"AB",X"65",X"A9",X"96",X"6A",X"A9",X"AA",
		X"AA",X"AE",X"FA",X"AA",X"AF",X"FE",X"EA",X"EF",
		X"AF",X"FE",X"EA",X"AB",X"BA",X"AA",X"AA",X"AA",
		X"AA",X"FE",X"BA",X"BA",X"AA",X"7A",X"AA",X"EB",
		X"EA",X"AF",X"AE",X"FA",X"AB",X"AB",X"6A",X"6A",
		X"A5",X"A5",X"59",X"55",X"A5",X"5A",X"AA",X"AA",
		X"9D",X"96",X"A5",X"59",X"96",X"A5",X"99",X"AA",
		X"AA",X"AA",X"AE",X"EA",X"FE",X"AA",X"B9",X"9A",
		X"EB",X"AA",X"AA",X"FE",X"AA",X"AF",X"EA",X"EA",
		X"AA",X"AB",X"AA",X"AA",X"E6",X"75",X"9A",X"D7",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"66",X"65",
		X"A6",X"56",X"59",X"96",X"66",X"6A",X"96",X"69",
		X"59",X"AA",X"65",X"59",X"56",X"65",X"A9",X"EA",
		X"AA",X"EA",X"AB",X"AA",X"AA",X"97",X"B8",X"9E",
		X"E6",X"E9",X"AA",X"AA",X"FE",X"AE",X"EE",X"AA",
		X"AE",X"A6",X"A6",X"BF",X"A6",X"75",X"9E",X"93",
		X"AA",X"5A",X"95",X"AA",X"AA",X"9A",X"6A",X"66",
		X"56",X"65",X"A9",X"9A",X"55",X"A9",X"AA",X"AA",
		X"AE",X"96",X"6A",X"59",X"9A",X"55",X"69",X"95",
		X"9A",X"AA",X"9A",X"A6",X"FA",X"EA",X"35",X"5E",
		X"A7",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"AA",X"AF",X"9A",X"FE",X"AF",X"EA",X"EA",X"AE",
		X"AA",X"AA",X"AA",X"AF",X"39",X"5D",X"AB",X"AA",
		X"6A",X"5A",X"AA",X"59",X"69",X"65",X"69",X"A6",
		X"66",X"55",X"56",X"AA",X"59",X"AA",X"75",X"A9",
		X"97",X"A9",X"59",X"A6",X"A5",X"5A",X"6A",X"A5",
		X"69",X"6A",X"95",X"A9",X"BF",X"AA",X"9E",X"EB",
		X"BF",X"AE",X"AA",X"AA",X"EE",X"AB",X"BA",X"9A",
		X"9A",X"AA",X"AA",X"BF",X"FA",X"AB",X"AA",X"6A",
		X"59",X"A9",X"AA",X"A6",X"9A",X"A5",X"55",X"95",
		X"55",X"59",X"95",X"A5",X"5A",X"AA",X"AA",X"5A",
		X"9A",X"65",X"59",X"96",X"66",X"59",X"AA",X"95",
		X"AA",X"AA",X"66",X"66",X"AA",X"FA",X"AB",X"BE",
		X"AA",X"55",X"AA",X"AA",X"AA",X"AB",X"7A",X"AA",
		X"EA",X"AA",X"A5",X"9A",X"AA",X"AA",X"5A",X"95",
		X"A6",X"AA",X"66",X"6A",X"6A",X"55",X"65",X"56",
		X"A5",X"55",X"9A",X"65",X"A9",X"96",X"A9",X"5E",
		X"9A",X"69",X"69",X"96",X"65",X"59",X"95",X"6A",
		X"65",X"56",X"AA",X"A9",X"AA",X"96",X"6A",X"5A",
		X"A9",X"A5",X"AA",X"BF",X"AA",X"A7",X"69",X"6A",
		X"A9",X"AA",X"6A",X"A5",X"96",X"5A",X"95",X"AA",
		X"6A",X"AA",X"AA",X"A9",X"95",X"6A",X"59",X"95",
		X"55",X"59",X"95",X"95",X"5A",X"9A",X"7A",X"A9",
		X"A6",X"65",X"99",X"95",X"A6",X"5A",X"9A",X"55",
		X"AA",X"A9",X"56",X"AA",X"AA",X"A9",X"99",X"AA",
		X"AA",X"AA",X"AA",X"6A",X"AA",X"A6",X"A9",X"6E",
		X"99",X"AA",X"6A",X"59",X"56",X"A5",X"AA",X"AA",
		X"A9",X"95",X"6A",X"A5",X"9A",X"95",X"A9",X"56",
		X"A5",X"55",X"56",X"66",X"59",X"AA",X"7A",X"5A",
		X"9A",X"A5",X"59",X"AA",X"65",X"55",X"56",X"A5",
		X"6A",X"96",X"AA",X"AA",X"AE",X"AA",X"A6",X"6A",
		X"96",X"A5",X"AE",X"56",X"AA",X"A7",X"65",X"AA",
		X"BA",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"AA",X"50",X"14",X"85",X"61",X"69",X"AA",X"AA",
		X"AA",X"A6",X"9A",X"9A",X"55",X"55",X"55",X"55",
		X"59",X"95",X"95",X"5A",X"AA",X"A6",X"AA",X"96",
		X"A5",X"5A",X"96",X"65",X"A9",X"96",X"6A",X"A9",
		X"6A",X"AA",X"A9",X"AA",X"AA",X"61",X"08",X"45",
		X"51",X"A9",X"69",X"AA",X"67",X"39",X"5A",X"EE",
		X"5A",X"11",X"19",X"96",X"65",X"58",X"9A",X"6A",
		X"A9",X"AA",X"59",X"69",X"A5",X"59",X"56",X"66",
		X"55",X"5A",X"A5",X"6A",X"96",X"7A",X"99",X"9A",
		X"69",X"59",X"96",X"6A",X"55",X"AA",X"65",X"66",
		X"AA",X"AA",X"BA",X"6A",X"96",X"65",X"15",X"95",
		X"51",X"A9",X"65",X"9A",X"96",X"78",X"9A",X"AA",
		X"55",X"50",X"15",X"41",X"61",X"58",X"96",X"AA",
		X"9A",X"AA",X"AA",X"96",X"6A",X"65",X"96",X"55",
		X"59",X"99",X"55",X"59",X"AA",X"AA",X"5A",X"AA",
		X"A5",X"5A",X"AA",X"65",X"A9",X"96",X"A6",X"AA",
		X"AA",X"AA",X"AA",X"5A",X"86",X"61",X"15",X"41",
		X"51",X"E5",X"69",X"9A",X"A7",X"28",X"5E",X"A6",
		X"95",X"51",X"09",X"85",X"65",X"55",X"86",X"A5",
		X"A9",X"A6",X"6A",X"A6",X"56",X"59",X"55",X"66",
		X"55",X"96",X"66",X"A9",X"9A",X"A9",X"AA",X"A7",
		X"66",X"59",X"A6",X"66",X"A9",X"96",X"A9",X"AA",
		X"9A",X"AA",X"66",X"58",X"96",X"50",X"58",X"45",
		X"54",X"A5",X"28",X"9A",X"A7",X"28",X"8E",X"A6",
		X"56",X"54",X"04",X"85",X"65",X"18",X"86",X"66",
		X"66",X"56",X"66",X"6A",X"A5",X"55",X"9A",X"55",
		X"69",X"55",X"A9",X"55",X"AA",X"66",X"6A",X"AA",
		X"A9",X"A9",X"96",X"65",X"A5",X"9A",X"6A",X"59",
		X"AA",X"AA",X"65",X"14",X"56",X"51",X"05",X"55",
		X"51",X"E5",X"68",X"8E",X"A2",X"38",X"8A",X"A6",
		X"45",X"11",X"15",X"56",X"60",X"14",X"56",X"65",
		X"A9",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"A6",X"55",X"5A",X"65",X"65",X"95",X"55",X"55",
		X"56",X"66",X"59",X"AA",X"BA",X"AA",X"97",X"6A",
		X"99",X"9A",X"A9",X"99",X"96",X"95",X"A5",X"5A",
		X"AA",X"2A",X"14",X"96",X"51",X"58",X"41",X"51",
		X"A2",X"28",X"9A",X"A3",X"29",X"4E",X"A6",X"55",
		X"50",X"54",X"46",X"21",X"58",X"96",X"61",X"59",
		X"6A",X"A5",X"55",X"5A",X"55",X"56",X"65",X"65",
		X"96",X"6A",X"A9",X"9A",X"6A",X"6A",X"AA",X"A5",
		X"5A",X"AA",X"65",X"69",X"A6",X"66",X"5A",X"A9",
		X"9A",X"65",X"14",X"81",X"15",X"18",X"55",X"50",
		X"E1",X"68",X"8E",X"A2",X"38",X"8E",X"A6",X"55",
		X"11",X"15",X"81",X"51",X"18",X"81",X"61",X"69",
		X"95",X"55",X"99",X"95",X"59",X"59",X"65",X"55",
		X"5A",X"A5",X"99",X"9A",X"AA",X"AA",X"E6",X"6A",
		X"A9",X"96",X"6A",X"5A",X"99",X"99",X"A9",X"AA",
		X"56",X"65",X"58",X"85",X"55",X"54",X"46",X"91",
		X"A2",X"28",X"8E",X"A2",X"29",X"8E",X"66",X"51",
		X"11",X"18",X"55",X"60",X"15",X"86",X"51",X"98",
		X"96",X"6A",X"55",X"55",X"55",X"95",X"95",X"56",
		X"56",X"66",X"66",X"AA",X"6A",X"A9",X"AA",X"65",
		X"6A",X"A6",X"66",X"55",X"A6",X"A6",X"AA",X"AA",
		X"9A",X"61",X"04",X"85",X"11",X"15",X"41",X"55",
		X"A1",X"39",X"8E",X"96",X"28",X"8E",X"A7",X"45",
		X"55",X"04",X"85",X"55",X"04",X"86",X"65",X"58",
		X"6A",X"A9",X"55",X"66",X"65",X"95",X"95",X"59",
		X"AA",X"A5",X"6A",X"AA",X"A9",X"AA",X"AB",X"A9",
		X"A9",X"96",X"65",X"A9",X"96",X"6A",X"A9",X"AA",
		X"56",X"60",X"58",X"42",X"55",X"44",X"46",X"51",
		X"E1",X"68",X"8E",X"A2",X"28",X"8E",X"A2",X"51",
		X"11",X"15",X"55",X"11",X"58",X"85",X"50",X"58",
		X"AA",X"55",X"99",X"6A",X"55",X"59",X"65",X"65",
		X"66",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"66",X"A9",X"AB",X"AA",X"99",X"AA",X"6A",X"A9",
		X"A6",X"66",X"56",X"5A",X"A9",X"A5",X"AA",X"86",
		X"61",X"15",X"46",X"61",X"15",X"41",X"55",X"A1",
		X"38",X"8E",X"56",X"68",X"8E",X"A7",X"45",X"61",
		X"44",X"46",X"50",X"19",X"82",X"65",X"58",X"AA",
		X"69",X"65",X"56",X"69",X"A5",X"95",X"5A",X"99",
		X"A9",X"A9",X"9A",X"AA",X"6A",X"AB",X"BA",X"AA",
		X"96",X"AA",X"59",X"AA",X"A5",X"AA",X"AA",X"46",
		X"61",X"58",X"41",X"15",X"14",X"55",X"90",X"A2",
		X"38",X"9A",X"92",X"28",X"8E",X"A2",X"42",X"15",
		X"14",X"55",X"21",X"14",X"85",X"11",X"58",X"AA",
		X"AA",X"5A",X"A5",X"55",X"56",X"A6",X"56",X"9A",
		X"AA",X"69",X"AA",X"A9",X"AA",X"AA",X"A5",X"9A",
		X"9A",X"A9",X"59",X"95",X"AA",X"AA",X"6B",X"86",
		X"15",X"58",X"85",X"50",X"15",X"81",X"81",X"A2",
		X"38",X"8E",X"65",X"28",X"8A",X"A7",X"45",X"11",
		X"15",X"46",X"54",X"58",X"56",X"61",X"58",X"AA",
		X"A9",X"56",X"66",X"56",X"99",X"95",X"99",X"AA",
		X"66",X"AA",X"9A",X"66",X"99",X"EA",X"AA",X"AE",
		X"AA",X"A9",X"AA",X"96",X"AA",X"AA",X"5A",X"56",
		X"61",X"14",X"56",X"51",X"44",X"45",X"55",X"A1",
		X"78",X"8A",X"56",X"68",X"8E",X"A3",X"85",X"55",
		X"54",X"41",X"61",X"14",X"46",X"60",X"98",X"AA",
		X"A9",X"5A",X"A5",X"65",X"56",X"6A",X"69",X"A5",
		X"A6",X"6A",X"AA",X"AA",X"6A",X"AA",X"AA",X"AE",
		X"9A",X"BA",X"AA",X"AA",X"AA",X"AA",X"6A",X"86",
		X"55",X"58",X"45",X"54",X"54",X"41",X"51",X"A2",
		X"38",X"8E",X"55",X"24",X"8A",X"A7",X"41",X"11",
		X"15",X"55",X"50",X"59",X"45",X"61",X"A9",X"AA",
		X"5A",X"A9",X"66",X"66",X"AA",X"A6",X"AA",X"9A",
		X"6A",X"A9",X"96",X"69",X"AA",X"EA",X"AA",X"AA",
		X"AB",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"AA",X"AA",X"AA",X"BA",X"FA",X"AB",X"86",X"25",
		X"54",X"46",X"15",X"14",X"55",X"81",X"A2",X"38",
		X"8A",X"56",X"28",X"8E",X"A6",X"45",X"55",X"44",
		X"45",X"60",X"54",X"46",X"60",X"A8",X"AA",X"AA",
		X"56",X"AA",X"59",X"66",X"66",X"6A",X"AA",X"AA",
		X"6A",X"AA",X"6A",X"A9",X"AA",X"AA",X"AE",X"AA",
		X"BA",X"AA",X"EA",X"AA",X"EA",X"AF",X"86",X"65",
		X"14",X"95",X"11",X"15",X"51",X"91",X"E2",X"7C",
		X"9A",X"51",X"29",X"8A",X"A3",X"42",X"51",X"15",
		X"55",X"61",X"05",X"85",X"65",X"A9",X"A6",X"A9",
		X"9A",X"A5",X"66",X"9A",X"AA",X"AA",X"9A",X"AA",
		X"AA",X"AA",X"6A",X"59",X"96",X"66",X"AA",X"EA",
		X"AA",X"AE",X"BA",X"BA",X"BA",X"BB",X"46",X"61",
		X"19",X"41",X"55",X"18",X"55",X"90",X"E2",X"38",
		X"9E",X"15",X"28",X"8E",X"A7",X"45",X"15",X"14",
		X"41",X"55",X"54",X"42",X"61",X"A9",X"AA",X"6A",
		X"AA",X"AA",X"A9",X"A6",X"AA",X"5A",X"AA",X"A6",
		X"6A",X"AA",X"65",X"99",X"95",X"A9",X"A9",X"96",
		X"BA",X"AA",X"EF",X"AA",X"AA",X"FF",X"96",X"61",
		X"15",X"85",X"55",X"44",X"45",X"91",X"E2",X"28",
		X"9E",X"51",X"15",X"8A",X"67",X"41",X"65",X"54",
		X"81",X"55",X"14",X"86",X"61",X"A9",X"AA",X"A9",
		X"9A",X"6A",X"AA",X"9A",X"AA",X"A9",X"AA",X"AA",
		X"AA",X"AA",X"65",X"59",X"9A",X"65",X"99",X"96",
		X"EA",X"EE",X"AA",X"FA",X"AB",X"FE",X"5A",X"51",
		X"19",X"51",X"51",X"15",X"55",X"51",X"E1",X"3C",
		X"4A",X"55",X"29",X"8A",X"57",X"45",X"11",X"15",
		X"45",X"15",X"58",X"81",X"A1",X"EA",X"AA",X"AA",
		X"56",X"AA",X"A9",X"9A",X"6A",X"6A",X"AA",X"A6",
		X"AA",X"AB",X"65",X"99",X"96",X"65",X"59",X"AA",
		X"BA",X"BB",X"EA",X"AE",X"BE",X"FA",X"9B",X"61",
		X"15",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"45",X"15",X"54",X"45",X"54",X"A1",X"78",X"8A",
		X"66",X"28",X"8A",X"56",X"45",X"55",X"44",X"55",
		X"51",X"04",X"96",X"A5",X"AE",X"AA",X"AA",X"AA",
		X"AA",X"A9",X"AA",X"AA",X"A9",X"AA",X"AA",X"AA",
		X"AA",X"69",X"59",X"56",X"A5",X"AA",X"AA",X"EA",
		X"EA",X"AB",X"BB",X"AB",X"EE",X"AA",X"51",X"19",
		X"51",X"61",X"05",X"55",X"51",X"A4",X"38",X"8F",
		X"56",X"28",X"9E",X"16",X"91",X"11",X"15",X"45",
		X"54",X"18",X"85",X"A5",X"AA",X"AA",X"A9",X"9A",
		X"AA",X"9A",X"9A",X"AA",X"AA",X"AA",X"AA",X"A9",
		X"AB",X"25",X"59",X"96",X"69",X"99",X"EA",X"BA",
		X"BE",X"FA",X"AB",X"FE",X"FE",X"AA",X"65",X"54",
		X"46",X"55",X"54",X"45",X"55",X"A0",X"78",X"8A",
		X"A6",X"38",X"9E",X"15",X"55",X"51",X"54",X"56",
		X"51",X"58",X"86",X"F5",X"AB",X"AB",X"AA",X"9A",
		X"AA",X"6A",X"AA",X"AA",X"A9",X"9A",X"AA",X"AA",
		X"AA",X"64",X"59",X"92",X"65",X"69",X"AA",X"AA",
		X"EA",X"AF",X"BE",X"AA",X"AA",X"AF",X"6A",X"18",
		X"55",X"61",X"55",X"81",X"55",X"A4",X"38",X"9A",
		X"A2",X"28",X"9A",X"06",X"56",X"51",X"19",X"55",
		X"60",X"54",X"86",X"AA",X"AA",X"AA",X"AA",X"A9",
		X"A6",X"AA",X"AB",X"A5",X"AA",X"A6",X"AA",X"AA",
		X"AB",X"65",X"49",X"A6",X"75",X"9A",X"9B",X"BA",
		X"BA",X"FA",X"AB",X"BF",X"AA",X"BB",X"66",X"15",
		X"56",X"61",X"15",X"55",X"51",X"A1",X"38",X"9A",
		X"62",X"38",X"9E",X"05",X"55",X"11",X"68",X"85",
		X"61",X"19",X"96",X"AA",X"AE",X"AA",X"6A",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"6A",X"AA",X"BA",X"AA",
		X"DA",X"25",X"59",X"96",X"B9",X"59",X"A6",X"AA",
		X"AF",X"AA",X"AA",X"AA",X"AF",X"AA",X"AA",X"19",
		X"96",X"55",X"59",X"45",X"55",X"A1",X"39",X"8E",
		X"A2",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"29",X"8E",X"55",X"56",X"61",X"59",X"95",X"51",
		X"59",X"9A",X"A5",X"AA",X"BA",X"AA",X"AA",X"AA",
		X"6A",X"AA",X"AA",X"A9",X"A6",X"A6",X"AE",X"AA",
		X"64",X"99",X"96",X"79",X"99",X"DA",X"EA",X"EA",
		X"EF",X"AE",X"AA",X"BA",X"AB",X"AA",X"59",X"96",
		X"66",X"68",X"45",X"95",X"E1",X"28",X"9A",X"A2",
		X"28",X"9A",X"56",X"56",X"61",X"69",X"96",X"55",
		X"68",X"96",X"A6",X"AA",X"EA",X"AA",X"AA",X"A6",
		X"AA",X"AA",X"A5",X"AA",X"9A",X"AA",X"AA",X"AA",
		X"64",X"49",X"97",X"64",X"59",X"EA",X"BE",X"AA",
		X"AA",X"BB",X"AA",X"EA",X"EA",X"6A",X"69",X"96",
		X"56",X"55",X"46",X"85",X"E2",X"28",X"8E",X"A2",
		X"28",X"8E",X"66",X"45",X"A5",X"15",X"85",X"A5",
		X"59",X"96",X"66",X"A9",X"9A",X"6A",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"AA",
		X"25",X"59",X"92",X"25",X"99",X"A6",X"AA",X"AA",
		X"AA",X"AA",X"A5",X"AA",X"AA",X"AA",X"59",X"9A",
		X"66",X"59",X"15",X"8A",X"E6",X"68",X"8A",X"A6",
		X"68",X"8A",X"97",X"85",X"65",X"55",X"9A",X"A5",
		X"59",X"9A",X"6A",X"A9",X"AA",X"AA",X"6A",X"A6",
		X"AA",X"EA",X"AA",X"99",X"AA",X"A5",X"AA",X"AA",
		X"64",X"49",X"96",X"64",X"99",X"9B",X"AA",X"AA",
		X"56",X"55",X"65",X"A9",X"AA",X"A6",X"AA",X"5A",
		X"9A",X"A2",X"28",X"8E",X"A3",X"38",X"8A",X"A2",
		X"28",X"8E",X"A2",X"68",X"56",X"19",X"9A",X"A5",
		X"A9",X"96",X"A6",X"99",X"AA",X"6A",X"66",X"66",
		X"6A",X"AA",X"AA",X"AA",X"AA",X"AA",X"99",X"9A",
		X"64",X"4C",X"92",X"60",X"99",X"96",X"BA",X"6A",
		X"56",X"55",X"59",X"A9",X"AB",X"6A",X"69",X"29",
		X"8A",X"A2",X"28",X"8A",X"A7",X"28",X"9A",X"A2",
		X"38",X"8A",X"A3",X"38",X"8A",X"A6",X"96",X"66",
		X"69",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"9A",X"6A",X"6A",X"96",X"A5",X"9A",X"5A",X"A9",
		X"A9",X"A6",X"AA",X"AB",X"6A",X"6A",X"AA",X"25",
		X"59",X"D2",X"25",X"59",X"A7",X"AA",X"5A",X"95",
		X"66",X"55",X"A9",X"AA",X"A9",X"A5",X"39",X"9A",
		X"A2",X"29",X"9A",X"A1",X"28",X"8A",X"A2",X"28",
		X"9A",X"91",X"58",X"89",X"A2",X"99",X"95",X"59",
		X"96",X"66",X"69",X"AA",X"AA",X"55",X"AA",X"95",
		X"9A",X"A9",X"AA",X"AA",X"AA",X"A9",X"A6",X"64",
		X"09",X"96",X"64",X"9D",X"AA",X"A6",X"5A",X"56",
		X"55",X"55",X"99",X"AA",X"A6",X"A6",X"28",X"8E",
		X"E6",X"69",X"4A",X"66",X"58",X"85",X"56",X"58",
		X"89",X"A6",X"39",X"8A",X"A2",X"78",X"A5",X"59",
		X"9A",X"A9",X"99",X"5A",X"65",X"6A",X"66",X"AA",
		X"6A",X"A6",X"5A",X"AA",X"A5",X"5A",X"9A",X"25",
		X"59",X"D2",X"24",X"59",X"E6",X"7A",X"AA",X"96",
		X"65",X"55",X"59",X"AA",X"AA",X"A6",X"38",X"8E",
		X"A2",X"69",X"9E",X"A2",X"28",X"95",X"91",X"68",
		X"9A",X"A6",X"68",X"8A",X"E2",X"68",X"AA",X"95",
		X"9A",X"AA",X"95",X"9A",X"99",X"59",X"95",X"A5",
		X"9A",X"A9",X"A6",X"9A",X"5A",X"A9",X"95",X"64",
		X"09",X"96",X"74",X"59",X"A6",X"66",X"59",X"56",
		X"55",X"59",X"55",X"AA",X"AA",X"A5",X"29",X"9A",
		X"A2",X"28",X"9A",X"A6",X"68",X"8A",X"A2",X"68",
		X"8E",X"A2",X"28",X"8A",X"E2",X"69",X"6A",X"69",
		X"A6",X"66",X"6A",X"AA",X"A5",X"95",X"56",X"55",
		X"99",X"AA",X"5A",X"6A",X"A5",X"5A",X"99",X"64",
		X"49",X"93",X"25",X"59",X"A7",X"BA",X"9A",X"96",
		X"69",X"59",X"69",X"95",X"A5",X"AA",X"28",X"8E",
		X"66",X"28",X"8A",X"E6",X"28",X"4A",X"A6",X"28",
		X"8A",X"A2",X"28",X"8E",X"E2",X"68",X"AA",X"A9",
		X"6A",X"A5",X"AA",X"6A",X"6A",X"55",X"56",X"A5",
		X"56",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"6A",X"A5",X"9A",X"5A",X"A9",X"95",X"25",X"59",
		X"96",X"64",X"4D",X"A6",X"65",X"59",X"AA",X"65",
		X"55",X"55",X"95",X"AA",X"A6",X"29",X"8A",X"E2",
		X"28",X"8A",X"A2",X"29",X"9A",X"A1",X"28",X"9A",
		X"A2",X"28",X"8E",X"A3",X"69",X"6A",X"A9",X"AA",
		X"56",X"A9",X"95",X"55",X"95",X"55",X"55",X"55",
		X"A6",X"AA",X"66",X"66",X"65",X"66",X"15",X"59",
		X"92",X"25",X"59",X"A7",X"76",X"5A",X"96",X"64",
		X"55",X"56",X"56",X"55",X"69",X"29",X"8E",X"E2",
		X"68",X"8E",X"E2",X"28",X"8A",X"E2",X"28",X"8A",
		X"A2",X"38",X"8A",X"A3",X"A9",X"A5",X"AA",X"95",
		X"5A",X"55",X"99",X"99",X"55",X"56",X"55",X"5A",
		X"69",X"6A",X"66",X"66",X"6A",X"95",X"65",X"09",
		X"96",X"25",X"59",X"A6",X"65",X"6A",X"96",X"65",
		X"5A",X"55",X"59",X"55",X"99",X"59",X"9A",X"B2",
		X"38",X"CA",X"E3",X"29",X"8A",X"A3",X"39",X"8A",
		X"A3",X"29",X"8E",X"A6",X"A9",X"95",X"A9",X"56",
		X"95",X"55",X"A6",X"5A",X"55",X"55",X"59",X"95",
		X"A6",X"AA",X"96",X"56",X"6A",X"55",X"64",X"55",
		X"95",X"64",X"5A",X"97",X"75",X"59",X"E6",X"69",
		X"55",X"56",X"55",X"55",X"55",X"55",X"85",X"A6",
		X"28",X"8E",X"E2",X"68",X"8A",X"A2",X"38",X"8E",
		X"E2",X"28",X"9E",X"A6",X"5A",X"69",X"55",X"69",
		X"55",X"6A",X"95",X"55",X"55",X"65",X"55",X"56",
		X"A5",X"56",X"AA",X"6A",X"69",X"95",X"55",X"49",
		X"96",X"25",X"59",X"92",X"69",X"99",X"AA",X"65",
		X"59",X"95",X"95",X"55",X"55",X"55",X"55",X"A5",
		X"29",X"9A",X"A2",X"29",X"8A",X"E2",X"28",X"8F",
		X"A2",X"68",X"9A",X"56",X"6A",X"55",X"55",X"95",
		X"5A",X"A9",X"55",X"55",X"59",X"65",X"55",X"A6",
		X"A5",X"99",X"5A",X"A5",X"56",X"6A",X"61",X"55",
		X"95",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"65",X"59",X"E6",X"65",X"5A",X"96",X"69",X"59",
		X"55",X"55",X"65",X"55",X"55",X"55",X"55",X"55",
		X"9A",X"A6",X"59",X"9A",X"A6",X"29",X"9A",X"A2",
		X"69",X"5A",X"55",X"55",X"55",X"55",X"95",X"A6",
		X"56",X"99",X"55",X"56",X"65",X"5A",X"9A",X"6A",
		X"A5",X"AA",X"95",X"99",X"99",X"55",X"55",X"56",
		X"65",X"49",X"96",X"65",X"99",X"96",X"65",X"5A",
		X"A5",X"55",X"5A",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"56",
		X"55",X"55",X"55",X"54",X"55",X"A5",X"55",X"A9",
		X"59",X"55",X"55",X"59",X"65",X"A5",X"96",X"A9",
		X"5A",X"5A",X"6A",X"65",X"56",X"65",X"55",X"95",
		X"55",X"99",X"96",X"65",X"5A",X"96",X"6A",X"5A",
		X"95",X"55",X"55",X"55",X"5A",X"59",X"55",X"58",
		X"55",X"51",X"55",X"55",X"55",X"54",X"55",X"65",
		X"55",X"45",X"55",X"55",X"5A",X"A9",X"95",X"56",
		X"99",X"95",X"5A",X"95",X"A9",X"99",X"96",X"AA",
		X"A9",X"AA",X"A5",X"66",X"6A",X"55",X"55",X"56",
		X"65",X"59",X"5A",X"65",X"A9",X"D6",X"69",X"A5",
		X"A6",X"55",X"59",X"55",X"55",X"55",X"55",X"65",
		X"8A",X"A6",X"68",X"8A",X"56",X"68",X"4A",X"A2",
		X"64",X"9A",X"56",X"59",X"A9",X"95",X"6A",X"A5",
		X"56",X"55",X"59",X"95",X"56",X"A9",X"AA",X"A9",
		X"95",X"5A",X"A9",X"95",X"99",X"A5",X"55",X"95",
		X"55",X"59",X"55",X"65",X"5A",X"9A",X"A9",X"99",
		X"96",X"65",X"55",X"45",X"55",X"55",X"55",X"55",
		X"95",X"A6",X"68",X"8A",X"92",X"68",X"8A",X"55",
		X"69",X"9A",X"56",X"95",X"9A",X"56",X"AA",X"55",
		X"55",X"6A",X"55",X"AA",X"A9",X"99",X"96",X"6A",
		X"A9",X"AA",X"95",X"6A",X"6A",X"55",X"66",X"66",
		X"65",X"55",X"99",X"95",X"99",X"A5",X"66",X"AA",
		X"A6",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"65",X"59",X"55",X"55",X"55",X"55",X"55",X"5A",
		X"A2",X"29",X"9A",X"A6",X"29",X"99",X"96",X"69",
		X"95",X"56",X"99",X"59",X"55",X"55",X"55",X"AA",
		X"A5",X"5A",X"96",X"6A",X"6A",X"AA",X"AA",X"5A",
		X"6A",X"66",X"AA",X"95",X"96",X"59",X"99",X"95",
		X"99",X"59",X"65",X"56",X"9A",X"A9",X"6A",X"EA",
		X"69",X"55",X"56",X"15",X"54",X"55",X"15",X"55",
		X"A5",X"55",X"49",X"A5",X"55",X"5A",X"55",X"59",
		X"55",X"99",X"55",X"56",X"55",X"55",X"5A",X"55",
		X"65",X"AA",X"9A",X"A9",X"A9",X"AA",X"6A",X"6A",
		X"A5",X"AA",X"AA",X"AA",X"95",X"56",X"55",X"56",
		X"55",X"59",X"99",X"59",X"A9",X"A5",X"9A",X"AA",
		X"6A",X"59",X"52",X"55",X"55",X"41",X"55",X"55",
		X"51",X"55",X"55",X"55",X"14",X"55",X"91",X"15",
		X"55",X"55",X"55",X"55",X"55",X"55",X"59",X"AA",
		X"A5",X"A9",X"A7",X"AA",X"9A",X"9A",X"AA",X"6A",
		X"AA",X"AA",X"A9",X"AA",X"AA",X"A5",X"9A",X"99",
		X"6A",X"55",X"A6",X"56",X"AA",X"AA",X"AD",X"AA",
		X"B9",X"9A",X"96",X"65",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"56",X"55",X"59",X"55",X"55",
		X"55",X"56",X"55",X"59",X"95",X"65",X"59",X"AA",
		X"B9",X"AA",X"EA",X"BA",X"AA",X"AB",X"AA",X"9A",
		X"AA",X"AA",X"AA",X"AA",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"FF",X"FF",X"FF",X"EA",X"AF",X"FA",X"AA",X"FE",
		X"EA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AB",
		X"6A",X"9A",X"A6",X"65",X"9A",X"9A",X"A9",X"9A",
		X"AA",X"A9",X"AA",X"EA",X"EF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"6A",X"9A",X"96",
		X"69",X"59",X"A6",X"A5",X"5A",X"A6",X"65",X"5A",
		X"AA",X"A9",X"9A",X"AA",X"A9",X"AA",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"AF",X"A6",X"65",X"5A",X"A6",
		X"55",X"5A",X"A6",X"65",X"9A",X"96",X"6A",X"9A",
		X"AA",X"B9",X"9A",X"AB",X"BA",X"AE",X"EA",X"EA",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"6A",X"5A",X"A6",X"65",X"5A",X"A6",
		X"65",X"5A",X"A6",X"65",X"5A",X"A6",X"69",X"99",
		X"96",X"A9",X"9E",X"EA",X"69",X"AA",X"EA",X"AE",
		X"AE",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AF",X"A6",X"65",X"5A",X"A2",X"65",X"9A",X"96",
		X"65",X"5A",X"96",X"59",X"99",X"96",X"69",X"99",
		X"A6",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"66",X"9A",X"EA",X"A9",X"AE",X"E6",X"AA",X"AE",
		X"FA",X"EB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"9A",
		X"96",X"25",X"59",X"A6",X"65",X"49",X"96",X"68",
		X"89",X"95",X"65",X"5A",X"96",X"65",X"5A",X"96",
		X"69",X"9E",X"96",X"6A",X"9A",X"AA",X"A9",X"AA",
		X"AB",X"BA",X"EA",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"25",X"59",
		X"52",X"54",X"49",X"92",X"25",X"5A",X"A6",X"65",
		X"49",X"A6",X"64",X"49",X"A5",X"65",X"5A",X"A6",
		X"65",X"99",X"A6",X"A5",X"5A",X"EA",X"A9",X"9A",
		X"EA",X"AA",X"AE",X"FA",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"EF",X"96",X"15",X"45",
		X"96",X"24",X"59",X"91",X"69",X"99",X"52",X"64",
		X"99",X"96",X"25",X"99",X"96",X"65",X"99",X"96",
		X"69",X"5A",X"EA",X"69",X"9E",X"A6",X"6A",X"AE",
		X"E6",X"AA",X"AF",X"EA",X"EA",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"5F",X"52",X"24",X"49",
		X"91",X"25",X"45",X"A6",X"24",X"59",X"A2",X"25",
		X"5A",X"92",X"69",X"49",X"A6",X"64",X"5A",X"A6",
		X"75",X"9A",X"E6",X"66",X"AA",X"EB",X"A9",X"AE",
		X"EA",X"AA",X"AE",X"FB",X"FA",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"49",X"91",X"25",X"59",
		X"96",X"24",X"59",X"92",X"64",X"49",X"92",X"69",
		X"99",X"92",X"25",X"55",X"96",X"79",X"5A",X"A6",
		X"69",X"9D",X"96",X"69",X"99",X"96",X"6A",X"AE",
		X"E6",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"A9",X"AE",X"EA",X"AE",X"AE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"25",X"45",X"96",X"14",X"45",X"51",
		X"14",X"45",X"51",X"15",X"45",X"52",X"25",X"49",
		X"56",X"64",X"49",X"55",X"65",X"49",X"96",X"69",
		X"99",X"96",X"69",X"99",X"96",X"A9",X"9A",X"AA",
		X"A9",X"AA",X"AB",X"BA",X"AE",X"FA",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"AB",X"14",X"44",X"41",X"14",X"04",X"51",
		X"10",X"05",X"41",X"10",X"05",X"51",X"10",X"05",
		X"51",X"14",X"45",X"91",X"14",X"55",X"52",X"65",
		X"55",X"96",X"65",X"59",X"A6",X"65",X"99",X"96",
		X"A9",X"9A",X"AA",X"AA",X"AA",X"AB",X"EA",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AF",X"42",X"10",X"05",X"41",X"10",X"05",X"41",
		X"10",X"44",X"41",X"14",X"04",X"51",X"10",X"45",
		X"41",X"54",X"44",X"45",X"54",X"59",X"55",X"64",
		X"45",X"66",X"65",X"56",X"96",X"A9",X"99",X"9A",
		X"A9",X"9A",X"EA",X"AA",X"AF",X"EA",X"EA",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"51",X"10",X"10",X"40",X"14",X"04",X"41",
		X"10",X"05",X"41",X"10",X"04",X"51",X"10",X"04",
		X"51",X"10",X"05",X"51",X"54",X"05",X"51",X"54",
		X"45",X"56",X"65",X"55",X"96",X"55",X"5A",X"A5",
		X"65",X"6A",X"A6",X"6A",X"AA",X"AA",X"AA",X"AA",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"51",X"10",X"10",X"50",X"10",X"10",X"50",
		X"40",X"40",X"01",X"01",X"44",X"41",X"14",X"44",
		X"41",X"14",X"55",X"41",X"54",X"05",X"95",X"10",
		X"55",X"56",X"25",X"55",X"95",X"54",X"99",X"95",
		X"69",X"95",X"9A",X"A9",X"9A",X"AA",X"A9",X"AA",
		X"EA",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"AA",X"AE",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"BF",X"4A",X"41",X"14",X"05",X"51",X"14",
		X"44",X"41",X"14",X"05",X"51",X"10",X"45",X"51",
		X"11",X"05",X"51",X"54",X"49",X"51",X"25",X"55",
		X"51",X"54",X"55",X"56",X"69",X"59",X"66",X"65",
		X"5A",X"AA",X"65",X"6A",X"A6",X"AA",X"9A",X"AB",
		X"AA",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"05",X"51",X"10",X"04",X"04",X"10",
		X"04",X"41",X"10",X"04",X"15",X"10",X"04",X"41",
		X"10",X"05",X"51",X"10",X"44",X"41",X"15",X"05",
		X"51",X"15",X"59",X"51",X"64",X"55",X"55",X"65",
		X"55",X"66",X"65",X"6A",X"A6",X"6A",X"AA",X"AA",
		X"AA",X"AF",X"EA",X"AA",X"FA",X"FF",X"FF",X"FF",
		X"FF",X"BF",X"4A",X"41",X"10",X"10",X"40",X"40",
		X"40",X"01",X"03",X"01",X"04",X"10",X"10",X"40",
		X"40",X"40",X"40",X"04",X"44",X"01",X"01",X"05",
		X"51",X"10",X"05",X"55",X"10",X"15",X"51",X"54",
		X"45",X"56",X"64",X"55",X"66",X"65",X"55",X"66",
		X"65",X"6A",X"A6",X"BA",X"AA",X"A6",X"AA",X"AA",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"9F",X"42",X"40",
		X"50",X"41",X"40",X"00",X"41",X"40",X"00",X"41",
		X"10",X"10",X"40",X"10",X"01",X"41",X"10",X"44",
		X"01",X"01",X"44",X"41",X"14",X"44",X"51",X"50",
		X"45",X"55",X"54",X"55",X"51",X"65",X"55",X"56",
		X"65",X"95",X"AA",X"A5",X"AA",X"A6",X"AA",X"9A",
		X"EA",X"AA",X"AE",X"AA",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"47",X"14",X"04",X"41",X"10",X"05",X"41",
		X"14",X"04",X"51",X"10",X"05",X"41",X"14",X"44",
		X"41",X"14",X"44",X"41",X"54",X"44",X"45",X"14",
		X"05",X"95",X"54",X"49",X"95",X"15",X"59",X"A5",
		X"55",X"5A",X"96",X"69",X"99",X"9A",X"A9",X"AA",
		X"AA",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"AA",X"AA",X"AB",X"EA",X"FF",X"FF",X"FF",X"AF",
		X"92",X"14",X"44",X"51",X"14",X"45",X"41",X"15",
		X"44",X"41",X"15",X"05",X"51",X"14",X"54",X"51",
		X"60",X"45",X"52",X"14",X"45",X"91",X"54",X"59",
		X"52",X"25",X"59",X"96",X"69",X"99",X"96",X"69",
		X"99",X"AA",X"AA",X"9A",X"AA",X"A9",X"AA",X"AB",
		X"7A",X"AB",X"AB",X"FA",X"FF",X"FF",X"FF",X"AF",
		X"92",X"25",X"49",X"91",X"64",X"49",X"96",X"24",
		X"05",X"52",X"14",X"48",X"95",X"24",X"05",X"52",
		X"25",X"44",X"52",X"21",X"59",X"52",X"25",X"49",
		X"96",X"65",X"99",X"96",X"69",X"5A",X"E6",X"69",
		X"AA",X"A6",X"79",X"AA",X"AB",X"7A",X"AE",X"EA",
		X"BE",X"AA",X"BB",X"BA",X"FB",X"FF",X"FF",X"9F",
		X"A7",X"39",X"49",X"96",X"14",X"49",X"92",X"69",
		X"99",X"53",X"20",X"55",X"92",X"65",X"49",X"92",
		X"24",X"5A",X"92",X"14",X"59",X"92",X"65",X"99",
		X"A6",X"68",X"5A",X"A2",X"65",X"9A",X"A7",X"7A",
		X"AE",X"A7",X"6A",X"AA",X"A7",X"BA",X"EA",X"FB",
		X"BA",X"AF",X"EB",X"BE",X"FE",X"FF",X"BF",X"9F",
		X"A7",X"78",X"5A",X"92",X"24",X"99",X"A6",X"34",
		X"9A",X"A7",X"65",X"9E",X"A2",X"79",X"9E",X"A6",
		X"65",X"9A",X"A7",X"79",X"4A",X"92",X"25",X"4A",
		X"96",X"79",X"99",X"A7",X"79",X"AA",X"A7",X"B9",
		X"AA",X"EB",X"B9",X"9E",X"EA",X"AE",X"EE",X"EB",
		X"BE",X"EE",X"BB",X"BB",X"FF",X"FF",X"BF",X"9B",
		X"E7",X"29",X"8D",X"E6",X"68",X"9D",X"93",X"68",
		X"49",X"E2",X"79",X"9A",X"E7",X"29",X"9A",X"E7",
		X"79",X"9E",X"E7",X"79",X"AE",X"E6",X"69",X"9A",
		X"E6",X"69",X"9E",X"D6",X"69",X"9E",X"EA",X"69",
		X"AE",X"E6",X"BA",X"AA",X"E7",X"BA",X"AF",X"FE",
		X"BA",X"BF",X"FB",X"BE",X"FA",X"FF",X"BF",X"9E",
		X"E6",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"24",X"5A",X"92",X"24",X"5A",X"A2",X"35",X"9A",
		X"93",X"29",X"49",X"92",X"10",X"54",X"A2",X"79",
		X"5E",X"A2",X"65",X"8A",X"E6",X"69",X"9E",X"A7",
		X"79",X"9A",X"A7",X"B9",X"99",X"A7",X"7A",X"9A",
		X"AB",X"BA",X"AF",X"FB",X"AA",X"EE",X"FB",X"BA",
		X"AB",X"AB",X"BA",X"EE",X"FF",X"7F",X"4A",X"92",
		X"24",X"49",X"92",X"24",X"49",X"92",X"24",X"49",
		X"92",X"24",X"49",X"41",X"10",X"44",X"95",X"24",
		X"59",X"92",X"25",X"59",X"92",X"64",X"59",X"96",
		X"65",X"99",X"96",X"69",X"5A",X"E6",X"65",X"AA",
		X"A6",X"69",X"AA",X"E6",X"BA",X"AA",X"AB",X"BA",
		X"AE",X"FA",X"BA",X"FA",X"FE",X"7F",X"49",X"96",
		X"20",X"05",X"41",X"14",X"44",X"92",X"14",X"48",
		X"91",X"14",X"49",X"41",X"14",X"45",X"92",X"25",
		X"49",X"91",X"24",X"45",X"52",X"15",X"49",X"95",
		X"64",X"5A",X"A6",X"65",X"9D",X"96",X"69",X"59",
		X"AA",X"B5",X"9A",X"AB",X"AA",X"AA",X"EA",X"AA",
		X"AA",X"AA",X"BE",X"AA",X"FF",X"7F",X"49",X"52",
		X"24",X"44",X"42",X"24",X"49",X"92",X"24",X"05",
		X"92",X"25",X"48",X"41",X"24",X"45",X"92",X"14",
		X"49",X"41",X"15",X"58",X"91",X"64",X"45",X"96",
		X"65",X"59",X"A6",X"65",X"9A",X"96",X"69",X"99",
		X"A6",X"6A",X"AA",X"A7",X"BA",X"AE",X"BB",X"BA",
		X"AA",X"EB",X"AA",X"EE",X"FE",X"7F",X"4A",X"92",
		X"14",X"09",X"91",X"24",X"49",X"52",X"20",X"49",
		X"91",X"24",X"49",X"92",X"15",X"49",X"96",X"24",
		X"55",X"92",X"14",X"09",X"91",X"15",X"59",X"96",
		X"69",X"89",X"97",X"69",X"9D",X"9A",X"79",X"AA",
		X"A7",X"7A",X"AE",X"EA",X"BA",X"AF",X"AB",X"BA",
		X"EE",X"FA",X"BA",X"AA",X"FF",X"7F",X"4A",X"96",
		X"24",X"59",X"92",X"24",X"49",X"96",X"24",X"59",
		X"92",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"24",X"49",X"92",X"24",X"45",X"96",X"64",X"49",
		X"96",X"64",X"59",X"92",X"65",X"9A",X"92",X"69",
		X"99",X"96",X"79",X"9A",X"E7",X"6A",X"AE",X"E6",
		X"BA",X"9A",X"EB",X"BE",X"EE",X"EB",X"BE",X"EE",
		X"EB",X"BE",X"EA",X"FF",X"7F",X"5A",X"A2",X"64",
		X"49",X"92",X"25",X"59",X"A2",X"25",X"4A",X"A6",
		X"64",X"49",X"96",X"64",X"49",X"A6",X"64",X"9E",
		X"A6",X"65",X"9A",X"E6",X"69",X"5E",X"E6",X"69",
		X"9E",X"A7",X"79",X"AA",X"AB",X"B9",X"9E",X"AB",
		X"B9",X"AE",X"FB",X"BA",X"AB",X"FB",X"BE",X"EA",
		X"EB",X"BE",X"FE",X"FF",X"7F",X"8A",X"97",X"29",
		X"9E",X"A2",X"64",X"4A",X"E6",X"24",X"99",X"93",
		X"29",X"5A",X"E6",X"68",X"8D",X"D6",X"39",X"5A",
		X"E3",X"29",X"9D",X"96",X"79",X"9A",X"E7",X"79",
		X"9E",X"EA",X"B9",X"9A",X"E7",X"6A",X"AE",X"EB",
		X"BE",X"EA",X"EB",X"BE",X"EE",X"EB",X"BE",X"FE",
		X"EB",X"AE",X"EE",X"FF",X"BF",X"4E",X"E6",X"64",
		X"4A",X"97",X"24",X"49",X"92",X"24",X"49",X"A2",
		X"25",X"9D",X"92",X"64",X"89",X"97",X"68",X"49",
		X"A6",X"64",X"5A",X"A3",X"79",X"9A",X"A7",X"B9",
		X"9A",X"A7",X"79",X"9A",X"AB",X"B9",X"9A",X"AB",
		X"B9",X"EE",X"EB",X"BA",X"AB",X"AB",X"BA",X"AB",
		X"FB",X"BA",X"BB",X"FF",X"BF",X"9A",X"E7",X"29",
		X"5E",X"A2",X"39",X"5A",X"A3",X"69",X"4E",X"E6",
		X"68",X"5E",X"E2",X"69",X"4A",X"E6",X"65",X"8E",
		X"D6",X"69",X"9E",X"E6",X"69",X"9E",X"A7",X"79",
		X"9A",X"EB",X"A9",X"9E",X"E6",X"6A",X"AE",X"FA",
		X"BA",X"AB",X"FB",X"BA",X"AE",X"FA",X"AA",X"AE",
		X"EA",X"AA",X"EF",X"FF",X"BF",X"AF",X"F7",X"79",
		X"9E",X"E7",X"79",X"EE",X"E7",X"79",X"EE",X"E7",
		X"7A",X"EF",X"EB",X"BD",X"EE",X"E7",X"7E",X"AF",
		X"FB",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"B9",X"EF",X"EB",X"BE",X"EE",X"EB",X"B9",X"AE",
		X"E7",X"BA",X"AF",X"FB",X"BA",X"EF",X"EB",X"BE",
		X"AF",X"FB",X"BE",X"AB",X"AB",X"BA",X"AE",X"EA",
		X"BF",X"FE",X"FF",X"FF",X"DF",X"AB",X"BD",X"DE",
		X"A7",X"69",X"9E",X"E6",X"69",X"9E",X"E6",X"7A",
		X"9A",X"F7",X"7A",X"9F",X"EA",X"69",X"9E",X"A6",
		X"79",X"9A",X"A7",X"79",X"9A",X"F7",X"BA",X"9B",
		X"FB",X"7A",X"EE",X"EB",X"BE",X"AF",X"FB",X"FE",
		X"EF",X"FF",X"BF",X"EE",X"EB",X"BE",X"EB",X"FB",
		X"FE",X"FF",X"FF",X"FF",X"AF",X"F7",X"79",X"9E",
		X"92",X"24",X"45",X"92",X"24",X"49",X"92",X"64",
		X"4A",X"96",X"64",X"99",X"E6",X"69",X"9D",X"E6",
		X"69",X"9E",X"E6",X"79",X"9F",X"AB",X"79",X"AA",
		X"E7",X"7A",X"AA",X"FB",X"B9",X"EA",X"FB",X"AA",
		X"EE",X"EB",X"BE",X"BF",X"FB",X"BF",X"FE",X"EF",
		X"BE",X"FE",X"FF",X"FF",X"AF",X"A6",X"B9",X"4A",
		X"52",X"10",X"49",X"95",X"14",X"55",X"A6",X"79",
		X"8A",X"96",X"68",X"49",X"A2",X"75",X"9A",X"E7",
		X"69",X"9E",X"A7",X"7A",X"9A",X"E6",X"69",X"9A",
		X"A6",X"B9",X"9A",X"A6",X"7A",X"AA",X"AB",X"BA",
		X"AF",X"EA",X"EE",X"EF",X"FB",X"BB",X"EF",X"FB",
		X"BB",X"FB",X"FF",X"FF",X"AF",X"A7",X"39",X"49",
		X"41",X"14",X"45",X"52",X"65",X"9E",X"E7",X"69",
		X"9E",X"E7",X"29",X"9E",X"92",X"79",X"9A",X"A7",
		X"B9",X"9E",X"E6",X"69",X"9E",X"E6",X"65",X"9E",
		X"E7",X"6A",X"AE",X"E7",X"6A",X"AE",X"FB",X"BA",
		X"AF",X"FF",X"BA",X"AF",X"AB",X"FE",X"EE",X"FF",
		X"FE",X"FF",X"FF",X"FF",X"EF",X"96",X"25",X"45",
		X"56",X"24",X"49",X"95",X"39",X"4A",X"92",X"24",
		X"89",X"E6",X"79",X"9E",X"E7",X"29",X"9D",X"96",
		X"69",X"5A",X"A7",X"65",X"5E",X"E6",X"6A",X"AE",
		X"EA",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"B9",X"EE",X"EA",X"BE",X"EE",X"EB",X"BE",X"EE",
		X"EB",X"FE",X"EE",X"FB",X"BF",X"EF",X"EB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"A7",X"24",X"55",X"92",
		X"54",X"49",X"A2",X"39",X"49",X"A2",X"24",X"49",
		X"92",X"69",X"9F",X"E7",X"79",X"9A",X"A7",X"79",
		X"9E",X"E6",X"79",X"AA",X"FB",X"B9",X"9E",X"FB",
		X"7A",X"AF",X"F7",X"BA",X"AF",X"FB",X"BE",X"EF",
		X"FA",X"BE",X"EF",X"FF",X"FA",X"EF",X"EF",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"EB",X"65",X"49",X"92",
		X"25",X"59",X"E6",X"24",X"59",X"A2",X"25",X"49",
		X"92",X"64",X"99",X"E6",X"7E",X"9E",X"E7",X"BE",
		X"EF",X"FB",X"BE",X"EF",X"EB",X"BE",X"EA",X"E7",
		X"6A",X"AA",X"AB",X"BE",X"EA",X"EB",X"EA",X"AF",
		X"FF",X"BB",X"FF",X"EB",X"BE",X"AF",X"FA",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"59",X"49",X"95",
		X"14",X"99",X"A3",X"74",X"8A",X"E7",X"78",X"9E",
		X"92",X"28",X"8D",X"A6",X"79",X"9A",X"AB",X"79",
		X"9A",X"A7",X"7A",X"9E",X"E6",X"69",X"9E",X"AA",
		X"A9",X"9E",X"AA",X"79",X"AA",X"AB",X"BA",X"AF",
		X"FB",X"AA",X"AF",X"BB",X"AA",X"AA",X"AB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"2A",X"45",X"51",
		X"54",X"59",X"A6",X"28",X"9D",X"E6",X"79",X"9E",
		X"93",X"25",X"5A",X"A7",X"79",X"89",X"A6",X"79",
		X"9A",X"E6",X"69",X"5A",X"A6",X"A9",X"9A",X"E7",
		X"6A",X"AE",X"E6",X"AA",X"AE",X"FA",X"BA",X"AA",
		X"BB",X"BA",X"AA",X"EA",X"BA",X"EA",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"19",X"95",
		X"10",X"45",X"91",X"69",X"9E",X"A7",X"78",X"9A",
		X"A7",X"64",X"9E",X"92",X"69",X"5A",X"A7",X"65",
		X"59",X"96",X"69",X"99",X"96",X"69",X"A9",X"96",
		X"A9",X"9A",X"AA",X"B9",X"EA",X"EB",X"BA",X"AB",
		X"AB",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"BA",X"EE",X"AB",X"BA",X"AA",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"BF",X"5B",X"52",X"65",
		X"49",X"91",X"64",X"89",X"E6",X"79",X"9E",X"E7",
		X"29",X"59",X"A6",X"64",X"99",X"96",X"65",X"5A",
		X"A6",X"65",X"99",X"96",X"6A",X"99",X"A6",X"6A",
		X"AE",X"AA",X"6A",X"AE",X"FA",X"AA",X"AE",X"EA",
		X"AA",X"AA",X"AB",X"BA",X"FB",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"96",X"29",
		X"59",X"56",X"25",X"5A",X"92",X"29",X"5A",X"A2",
		X"64",X"49",X"96",X"25",X"55",X"52",X"65",X"55",
		X"56",X"65",X"5A",X"A6",X"65",X"AA",X"96",X"6A",
		X"A9",X"A6",X"BA",X"AA",X"EA",X"BE",X"EE",X"EA",
		X"BE",X"AF",X"FA",X"FA",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A7",X"65",
		X"5A",X"A6",X"64",X"99",X"96",X"64",X"49",X"56",
		X"25",X"56",X"56",X"68",X"55",X"66",X"65",X"9A",
		X"96",X"A9",X"95",X"9A",X"69",X"A9",X"A6",X"AA",
		X"9E",X"EA",X"AA",X"AE",X"FA",X"AA",X"AF",X"AB",
		X"BA",X"AF",X"BB",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"69",
		X"99",X"96",X"69",X"49",X"56",X"65",X"5A",X"A2",
		X"65",X"99",X"95",X"65",X"5A",X"A6",X"55",X"99",
		X"95",X"69",X"5A",X"A6",X"A9",X"9A",X"EA",X"A9",
		X"AA",X"A6",X"BA",X"AA",X"AA",X"BA",X"EE",X"EA",
		X"FE",X"EA",X"EB",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"6A",
		X"5A",X"A6",X"65",X"5A",X"91",X"55",X"5A",X"A6",
		X"65",X"5A",X"A6",X"65",X"5A",X"A6",X"69",X"6A",
		X"A6",X"6A",X"A9",X"AA",X"6A",X"AA",X"AA",X"BA",
		X"AA",X"EB",X"AA",X"9B",X"AB",X"BE",X"AA",X"FB",
		X"AA",X"EE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"9A",
		X"96",X"69",X"99",X"96",X"65",X"5A",X"A6",X"25",
		X"99",X"96",X"69",X"99",X"96",X"69",X"99",X"96",
		X"A9",X"9A",X"A6",X"76",X"AA",X"A7",X"7A",X"AA",
		X"BB",X"BA",X"AE",X"EA",X"AA",X"AF",X"AB",X"BE",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"97",X"69",X"5A",X"A6",X"69",X"9A",X"A6",X"A9",
		X"5A",X"A6",X"69",X"9A",X"AA",X"BA",X"9A",X"AA",
		X"B9",X"9A",X"AB",X"BA",X"AA",X"EB",X"AA",X"AF",
		X"AB",X"BE",X"EE",X"AB",X"BE",X"FE",X"EB",X"FE",
		X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"6A",X"AA",X"A7",X"65",X"AA",X"EB",X"75",
		X"AA",X"A7",X"A9",X"99",X"EA",X"69",X"AA",X"E7",
		X"6A",X"AE",X"EA",X"BE",X"AE",X"FA",X"BE",X"AA",
		X"FB",X"EA",X"AF",X"FB",X"AA",X"EE",X"AB",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"BA",X"9A",X"EA",X"A9",X"9E",X"A6",X"6A",
		X"AE",X"EA",X"B9",X"9E",X"AB",X"B9",X"AA",X"AB",
		X"BA",X"AA",X"EB",X"AA",X"AF",X"EB",X"BE",X"BF",
		X"FB",X"BA",X"BF",X"EA",X"BF",X"FE",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"AF",X"AB",X"A9",X"5A",X"EA",X"A9",
		X"9E",X"E6",X"AA",X"9A",X"AA",X"7A",X"AA",X"E6",
		X"6A",X"AE",X"EA",X"BE",X"AA",X"BB",X"BA",X"AA",
		X"AB",X"BA",X"EA",X"EB",X"AA",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"FF",X"FF",X"EB",X"6A",X"AA",X"A6",X"66",X"AA",
		X"A6",X"66",X"AE",X"A6",X"6A",X"AA",X"AB",X"AA",
		X"AE",X"A6",X"BA",X"EA",X"AB",X"BA",X"AF",X"FA",
		X"BA",X"AB",X"BB",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"BF",X"AE",X"E6",X"6A",X"A9",
		X"E6",X"6A",X"6A",X"AA",X"B9",X"AA",X"A6",X"BA",
		X"EA",X"AB",X"BA",X"AF",X"EA",X"AA",X"AB",X"FB",
		X"AB",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AA",X"AE",
		X"AA",X"BA",X"AE",X"AB",X"BA",X"AE",X"EA",X"AA",
		X"AF",X"EA",X"BE",X"EA",X"EB",X"FE",X"AE",X"FE",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",
		X"FB",X"AA",X"AB",X"FB",X"AA",X"AF",X"FB",X"BE",
		X"EE",X"FB",X"AB",X"AF",X"FF",X"EA",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"BF",X"FA",X"AF",X"FE",X"EA",
		X"AF",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"18",X"00",X"FB",X"EE",X"19",X"02",X"00",
		X"E5",X"1A",X"21",X"E6",X"20",X"35",X"53",X"0B",
		X"21",X"0E",X"F3",X"17",X"90",X"05",X"59",X"00",
		X"2B",X"30",X"CD",X"5F",X"21",X"32",X"E6",X"52",
		X"35",X"53",X"21",X"E3",X"32",X"2B",X"34",X"11",
		X"00",X"07",X"90",X"26",X"2B",X"34",X"11",X"00",
		X"08",X"2B",X"36",X"21",X"34",X"E9",X"E9",X"99",
		X"34",X"99",X"36",X"2B",X"36",X"21",X"38",X"5E",
		X"24",X"21",X"3A",X"5E",X"25",X"21",X"3C",X"2B",
		X"28",X"E3",X"06",X"2B",X"3C",X"11",X"E1",X"04",
		X"2B",X"22",X"59",X"FB",X"2B",X"34",X"21",X"36",
		X"7F",X"00",X"93",X"36",X"5E",X"26",X"B4",X"CB",
		X"93",X"28",X"93",X"34",X"21",X"34",X"35",X"72",
		X"4B",X"FF",X"2B",X"3E",X"CD",X"76",X"75",X"2B",
		X"40",X"21",X"40",X"AD",X"2B",X"32",X"93",X"40",
		X"35",X"3F",X"74",X"CF",X"3E",X"90",X"66",X"63",
		X"FF",X"2B",X"42",X"CD",X"90",X"35",X"56",X"8F",
		X"2B",X"34",X"21",X"3A",X"F0",X"3C",X"21",X"3C",
		X"99",X"44",X"2B",X"3C",X"21",X"34",X"E6",X"01",
		X"90",X"7A",X"FF",X"2B",X"46",X"CD",X"BC",X"75",
		X"1A",X"0E",X"B8",X"48",X"82",X"80",X"35",X"72",
		X"A9",X"21",X"4A",X"35",X"56",X"A7",X"E6",X"01",
		X"2B",X"4A",X"CF",X"4C",X"1A",X"11",X"82",X"80",
		X"35",X"72",X"B4",X"E6",X"01",X"90",X"B6",X"59",
		X"00",X"99",X"4E",X"CF",X"50",X"63",X"FF",X"2B",
		X"52",X"CD",X"DE",X"75",X"11",X"20",X"08",X"2B",
		X"3C",X"59",X"08",X"2B",X"3A",X"59",X"00",X"2B",
		X"38",X"21",X"4A",X"2B",X"54",X"CF",X"56",X"21",
		X"48",X"E3",X"3C",X"82",X"FF",X"2B",X"48",X"63",
		X"FF",X"2B",X"4C",X"93",X"1B",X"FF",X"03",X"00",
		X"F7",X"CD",X"0B",X"00",X"FD",X"04",X"68",X"18",
		X"75",X"59",X"0F",X"2B",X"3A",X"21",X"58",X"CF",
		X"5A",X"63",X"FF",X"2B",X"5C",X"CD",X"43",X"75",
		X"11",X"35",X"44",X"2B",X"3C",X"59",X"04",X"2B",
		X"38",X"CD",X"25",X"47",X"41",X"4D",X"45",X"20",
		X"4F",X"56",X"45",X"52",X"00",X"CF",X"42",X"21",
		X"5E",X"B8",X"30",X"35",X"56",X"3F",X"21",X"60",
		X"FC",X"62",X"35",X"72",X"3F",X"21",X"5E",X"2B",
		X"30",X"59",X"1E",X"2B",X"3A",X"CF",X"64",X"CF",
		X"66",X"63",X"FF",X"2B",X"68",X"CD",X"59",X"2B",
		X"6A",X"1A",X"0E",X"99",X"6A",X"82",X"FF",X"2B",
		X"6A",X"1A",X"0E",X"B8",X"6A",X"35",X"72",X"51",
		X"FF",X"2B",X"50",X"CD",X"7F",X"75",X"59",X"08",
		X"2B",X"3A",X"59",X"00",X"2B",X"38",X"11",X"00",
		X"08",X"CF",X"6C",X"11",X"38",X"08",X"2B",X"3C",
		X"CD",X"7B",X"47",X"69",X"67",X"61",X"74",X"72",
		X"6F",X"6E",X"00",X"CF",X"42",X"63",X"FF",X"2B",
		X"6E",X"CD",X"A3",X"2B",X"70",X"11",X"03",X"0B",
		X"2B",X"22",X"21",X"38",X"5E",X"25",X"21",X"70",
		X"2B",X"26",X"59",X"A0",X"5E",X"24",X"B4",X"F3",
		X"11",X"00",X"01",X"99",X"70",X"2B",X"70",X"35",
		X"4D",X"90",X"FF",X"2B",X"6C",X"CD",X"C1",X"59",
		X"00",X"B8",X"72",X"2B",X"6A",X"21",X"74",X"2B",
		X"72",X"21",X"6A",X"2B",X"74",X"21",X"76",X"35",
		X"53",X"BC",X"59",X"00",X"E3",X"3C",X"2B",X"76",
		X"FF",X"2B",X"78",X"CD",X"DF",X"59",X"00",X"B8",
		X"74",X"2B",X"6A",X"21",X"72",X"2B",X"74",X"21",
		X"6A",X"2B",X"72",X"21",X"76",X"35",X"56",X"DA",
		X"59",X"00",X"E6",X"3C",X"2B",X"76",X"FF",X"2B",
		X"7A",X"CD",X"F0",X"2B",X"3C",X"21",X"3A",X"5E",
		X"19",X"F3",X"3C",X"93",X"3D",X"F3",X"3C",X"FF",
		X"2B",X"5A",X"93",X"1B",X"FF",X"04",X"00",X"F9",
		X"CD",X"AE",X"75",X"00",X"FD",X"04",X"68",X"18",
		X"CF",X"60",X"1A",X"75",X"82",X"80",X"2B",X"6A",
		X"21",X"74",X"82",X"02",X"35",X"3F",X"12",X"59",
		X"40",X"99",X"6A",X"E3",X"1B",X"2B",X"3A",X"1A",
		X"59",X"FC",X"58",X"82",X"02",X"35",X"3F",X"23",
		X"59",X"01",X"FC",X"3A",X"2B",X"3A",X"21",X"58",
		X"CF",X"5A",X"21",X"58",X"99",X"74",X"2B",X"58",
		X"21",X"58",X"AD",X"82",X"03",X"35",X"3F",X"3B",
		X"63",X"FF",X"21",X"58",X"AD",X"8C",X"18",X"35",
		X"72",X"5D",X"59",X"40",X"99",X"4A",X"CF",X"7C",
		X"59",X"02",X"5E",X"2C",X"21",X"5E",X"99",X"4A",
		X"2B",X"5E",X"CF",X"7E",X"59",X"05",X"CF",X"81",
		X"93",X"83",X"93",X"85",X"CF",X"5C",X"21",X"83",
		X"35",X"56",X"6C",X"E6",X"01",X"2B",X"83",X"CF",
		X"87",X"90",X"AA",X"21",X"89",X"AD",X"2B",X"6A",
		X"21",X"85",X"35",X"56",X"7E",X"E6",X"01",X"2B",
		X"85",X"59",X"3E",X"90",X"80",X"59",X"04",X"2B",
		X"3A",X"21",X"89",X"CF",X"5A",X"21",X"6A",X"82",
		X"40",X"35",X"72",X"92",X"11",X"00",X"01",X"90",
		X"94",X"59",X"01",X"2B",X"8B",X"21",X"6A",X"82",
		X"80",X"35",X"72",X"A1",X"21",X"8B",X"90",X"A5",
		X"59",X"00",X"B8",X"8B",X"E9",X"99",X"89",X"2B",
		X"89",X"CF",X"52",X"90",X"01",X"2B",X"8D",X"CD",
		X"EE",X"75",X"59",X"18",X"2B",X"3A",X"11",X"A7",
		X"04",X"2B",X"22",X"B4",X"FD",X"2B",X"3C",X"1A",
		X"3C",X"E6",X"80",X"35",X"53",X"C9",X"E3",X"96",
		X"E3",X"05",X"82",X"FE",X"5E",X"3C",X"1A",X"3D",
		X"82",X"7F",X"E6",X"40",X"35",X"53",X"DA",X"E3",
		X"66",X"E3",X"15",X"82",X"FE",X"5E",X"3D",X"21",
		X"3C",X"AD",X"8C",X"04",X"35",X"72",X"B7",X"21",
		X"3C",X"CF",X"5A",X"63",X"FF",X"2B",X"87",X"59",
		X"00",X"2B",X"76",X"93",X"1B",X"FF",X"05",X"00",
		X"ED",X"CD",X"E6",X"00",X"FD",X"04",X"68",X"18",
		X"75",X"1A",X"11",X"82",X"CF",X"8C",X"CF",X"35",
		X"3F",X"0E",X"CF",X"8F",X"63",X"FF",X"21",X"78",
		X"2B",X"70",X"21",X"7A",X"2B",X"91",X"21",X"58",
		X"99",X"74",X"AD",X"8C",X"04",X"2B",X"6A",X"35",
		X"3F",X"2B",X"8C",X"1C",X"35",X"72",X"29",X"2B",
		X"6A",X"90",X"39",X"21",X"58",X"99",X"74",X"99",
		X"74",X"AD",X"8C",X"3E",X"35",X"72",X"39",X"93",
		X"6B",X"21",X"58",X"B8",X"72",X"AD",X"8C",X"04",
		X"35",X"3F",X"54",X"8C",X"1C",X"35",X"72",X"4E",
		X"2B",X"91",X"93",X"6B",X"90",X"52",X"59",X"00",
		X"2B",X"70",X"90",X"71",X"21",X"58",X"B8",X"72",
		X"B8",X"72",X"AD",X"8C",X"04",X"35",X"3F",X"71",
		X"8C",X"1C",X"35",X"72",X"6B",X"2B",X"91",X"93",
		X"6B",X"90",X"71",X"21",X"76",X"E3",X"0F",X"21",
		X"76",X"21",X"58",X"99",X"72",X"AD",X"8C",X"04",
		X"35",X"3F",X"8C",X"8C",X"1C",X"35",X"72",X"86",
		X"2B",X"70",X"93",X"6B",X"90",X"8A",X"59",X"00",
		X"2B",X"91",X"90",X"A9",X"21",X"58",X"99",X"72",
		X"99",X"72",X"AD",X"8C",X"04",X"35",X"3F",X"A9",
		X"8C",X"1C",X"35",X"72",X"A3",X"2B",X"70",X"93",
		X"6B",X"90",X"A9",X"21",X"76",X"E6",X"0F",X"21",
		X"76",X"21",X"6A",X"35",X"72",X"BB",X"1A",X"06",
		X"E6",X"0D",X"35",X"53",X"B9",X"59",X"01",X"90",
		X"BB",X"59",X"00",X"35",X"3F",X"E4",X"21",X"70",
		X"35",X"72",X"C7",X"21",X"91",X"90",X"DF",X"21",
		X"91",X"35",X"72",X"D0",X"21",X"70",X"90",X"DF",
		X"1A",X"06",X"E6",X"80",X"99",X"76",X"35",X"53",
		X"DD",X"21",X"70",X"90",X"DF",X"21",X"91",X"35",
		X"3F",X"E4",X"CF",X"18",X"63",X"FF",X"2B",X"93",
		X"93",X"1B",X"FF",X"06",X"00",X"FA",X"CD",X"16",
		X"75",X"99",X"4A",X"2B",X"4A",X"E6",X"0F",X"35",
		X"56",X"0E",X"59",X"00",X"FD",X"04",X"68",X"18",
		X"0F",X"2B",X"4A",X"1A",X"0E",X"2B",X"48",X"CF",
		X"4C",X"63",X"FF",X"2B",X"81",X"CD",X"B3",X"75",
		X"59",X"00",X"2B",X"5E",X"2B",X"4A",X"CF",X"7E",
		X"59",X"0F",X"2B",X"4A",X"CF",X"4C",X"CF",X"64",
		X"59",X"04",X"2B",X"38",X"11",X"00",X"10",X"2B",
		X"3C",X"CF",X"6C",X"59",X"1A",X"2B",X"3A",X"59",
		X"01",X"2B",X"44",X"59",X"9F",X"CF",X"46",X"11",
		X"00",X"01",X"2B",X"44",X"59",X"6F",X"CF",X"46",
		X"11",X"FF",X"FF",X"2B",X"44",X"59",X"9F",X"CF",
		X"46",X"11",X"00",X"FF",X"2B",X"44",X"59",X"6E",
		X"CF",X"46",X"59",X"01",X"2B",X"44",X"59",X"9E",
		X"CF",X"46",X"11",X"00",X"01",X"2B",X"44",X"59",
		X"6D",X"CF",X"46",X"11",X"FF",X"FF",X"2B",X"44",
		X"59",X"9D",X"CF",X"46",X"11",X"00",X"FF",X"2B",
		X"44",X"59",X"6D",X"CF",X"46",X"CF",X"95",X"11",
		X"30",X"44",X"2B",X"58",X"2B",X"89",X"CF",X"5C",
		X"59",X"00",X"2B",X"83",X"2B",X"85",X"2B",X"4A",
		X"59",X"0F",X"CF",X"81",X"59",X"02",X"2B",X"74",
		X"11",X"00",X"02",X"2B",X"72",X"59",X"19",X"2B",
		X"34",X"CF",X"87",X"21",X"34",X"E6",X"01",X"35",
		X"4D",X"A2",X"21",X"97",X"2B",X"60",X"63",X"FF",
		X"2B",X"8F",X"CD",X"F0",X"75",X"11",X"02",X"08",
		X"2B",X"3C",X"21",X"5E",X"B8",X"30",X"35",X"56",
		X"C8",X"59",X"1E",X"90",X"CA",X"59",X"08",X"2B",
		X"3A",X"59",X"00",X"2B",X"38",X"21",X"5E",X"2B",
		X"54",X"CF",X"99",X"21",X"5E",X"E6",X"64",X"35",
		X"53",X"E1",X"59",X"04",X"90",X"EC",X"E6",X"C8",
		X"35",X"53",X"EA",X"59",X"03",X"90",X"EC",X"59",
		X"02",X"2B",X"4E",X"63",X"FF",X"2B",X"7E",X"11",
		X"A0",X"08",X"2B",X"1A",X"FF",X"08",X"A0",X"56",
		X"CD",X"D4",X"75",X"11",X"9C",X"44",X"B8",X"58",
		X"35",X"72",X"C3",X"00",X"FD",X"04",X"68",X"18",
		X"59",X"1E",X"2B",X"3A",X"11",X"02",X"08",X"2B",
		X"3C",X"CD",X"B9",X"41",X"55",X"54",X"4F",X"00",
		X"CF",X"42",X"21",X"93",X"2B",X"60",X"CF",X"18",
		X"90",X"D2",X"1A",X"11",X"82",X"CF",X"8C",X"CF",
		X"35",X"3F",X"D2",X"21",X"62",X"2B",X"60",X"CF",
		X"18",X"63",X"FF",X"2B",X"97",X"CD",X"EF",X"75",
		X"59",X"20",X"2B",X"32",X"59",X"0A",X"2B",X"9B",
		X"CF",X"9D",X"59",X"30",X"2B",X"32",X"59",X"01",
		X"2B",X"9B",X"CF",X"9D",X"63",X"FF",X"2B",X"56",
		X"93",X"1B",X"FF",X"09",X"A0",X"56",X"CD",X"C7",
		X"75",X"21",X"54",X"B8",X"9B",X"35",X"50",X"C3",
		X"2B",X"54",X"59",X"31",X"2B",X"32",X"21",X"54",
		X"B8",X"9B",X"35",X"50",X"BB",X"2B",X"54",X"93",
		X"32",X"90",X"B0",X"CF",X"3E",X"59",X"30",X"2B",
		X"32",X"90",X"C5",X"CF",X"3E",X"63",X"FF",X"2B",
		X"9D",X"CD",X"EF",X"75",X"59",X"20",X"2B",X"32",
		X"11",X"E8",X"03",X"2B",X"9B",X"CF",X"9D",X"59",
		X"64",X"2B",X"9B",X"CF",X"9D",X"59",X"0A",X"2B",
		X"9B",X"CF",X"9D",X"59",X"30",X"2B",X"32",X"59",
		X"01",X"2B",X"9B",X"CF",X"9D",X"63",X"FF",X"2B",
		X"99",X"93",X"1B",X"FF",X"0A",X"A0",X"56",X"CD",
		X"BA",X"75",X"11",X"74",X"08",X"2B",X"3C",X"59",
		X"00",X"2B",X"38",X"CD",X"B0",X"48",X"49",X"20",
		X"00",X"CF",X"42",X"21",X"30",X"2B",X"54",X"CF",
		X"99",X"63",X"FF",X"2B",X"64",X"CD",X"EF",X"2B",
		X"34",X"88",X"FF",X"8C",X"FF",X"88",X"FA",X"2B",
		X"70",X"1A",X"34",X"2B",X"34",X"59",X"00",X"F0",
		X"70",X"93",X"70",X"59",X"01",X"F0",X"70",X"93",
		X"70",X"11",X"00",X"09",X"99",X"34",X"7F",X"00",
		X"F0",X"70",X"93",X"70",X"11",X"00",X"09",X"99",
		X"34",X"7F",X"01",X"F0",X"70",X"93",X"70",X"FF",
		X"2B",X"9F",X"93",X"00",X"FD",X"04",X"68",X"18",
		X"1B",X"FF",X"0B",X"A0",X"4C",X"CD",X"C2",X"75",
		X"E9",X"2B",X"6A",X"11",X"00",X"01",X"FA",X"6A",
		X"CF",X"9F",X"11",X"00",X"02",X"FA",X"6A",X"CF",
		X"9F",X"11",X"00",X"03",X"FA",X"6A",X"CF",X"9F",
		X"11",X"00",X"04",X"FA",X"6A",X"CF",X"9F",X"63",
		X"FF",X"2B",X"7C",X"CD",X"E5",X"75",X"59",X"49",
		X"2B",X"A1",X"21",X"A1",X"CF",X"7C",X"59",X"05",
		X"5E",X"2C",X"1A",X"2C",X"35",X"72",X"D3",X"21",
		X"A1",X"E6",X"01",X"2B",X"A1",X"8C",X"30",X"35",
		X"72",X"CB",X"63",X"FF",X"2B",X"66",X"93",X"1B",
		X"FF",X"0C",X"A0",X"45",X"CD",X"DE",X"75",X"11",
		X"33",X"45",X"2B",X"70",X"2B",X"3C",X"59",X"18",
		X"2B",X"3A",X"21",X"A3",X"CF",X"42",X"59",X"2D",
		X"CF",X"50",X"21",X"70",X"2B",X"3C",X"59",X"3E",
		X"2B",X"3A",X"21",X"40",X"CF",X"42",X"59",X"2D",
		X"CF",X"50",X"21",X"70",X"2B",X"3C",X"59",X"0F",
		X"2B",X"3A",X"21",X"40",X"CF",X"42",X"59",X"2D",
		X"CF",X"50",X"21",X"70",X"2B",X"3C",X"21",X"40",
		X"CF",X"42",X"63",X"FF",X"2B",X"95",X"93",X"1B",
		X"FF",X"0D",X"A0",X"46",X"CD",X"DF",X"21",X"74",
		X"2B",X"6A",X"1A",X"11",X"8C",X"FE",X"35",X"72",
		X"AF",X"59",X"02",X"2B",X"6A",X"1A",X"11",X"8C",
		X"FD",X"35",X"72",X"BB",X"11",X"FE",X"FF",X"2B",
		X"6A",X"1A",X"11",X"8C",X"FB",X"35",X"72",X"C7",
		X"11",X"00",X"02",X"2B",X"6A",X"1A",X"11",X"8C",
		X"F7",X"35",X"72",X"D3",X"11",X"00",X"FE",X"2B",
		X"6A",X"21",X"6A",X"99",X"74",X"35",X"3F",X"DE",
		X"21",X"6A",X"2B",X"74",X"FF",X"2B",X"62",X"93",
		X"1B",X"FF",X"0E",X"A0",X"4D",X"CD",X"CB",X"20",
		X"45",X"41",X"54",X"20",X"46",X"4F",X"4F",X"44",
		X"00",X"4E",X"4F",X"54",X"20",X"50",X"4F",X"49",
		X"53",X"4F",X"4E",X"00",X"FD",X"04",X"68",X"18",
		X"00",X"47",X"45",X"54",X"20",X"52",X"45",X"41",
		X"44",X"59",X"21",X"00",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"2B",
		X"A3",X"CF",X"6E",X"59",X"49",X"CF",X"7C",X"CF",
		X"8F",X"CF",X"8D",X"59",X"78",X"5E",X"2C",X"59",
		X"07",X"2B",X"3A",X"21",X"58",X"CF",X"5A",X"CF",
		X"68",X"59",X"3C",X"CF",X"50",X"90",X"D3",X"00",
		X"26",X"27",X"00",X"1D",X"28",X"24",X"25",X"00",
		X"24",X"04",X"24",X"1D",X"28",X"26",X"01",X"26",
		X"4C",X"16",X"4E",X"00",X"02",X"16",X"03",X"CB",
		X"EC",X"27",X"08",X"56",X"57",X"00",X"01",X"1D",
		X"25",X"24",X"02",X"24",X"EE",X"18",X"19",X"26",
		X"FE",X"1D",X"00",X"26",X"01",X"26",X"03",X"CB",
		X"EC",X"53",X"6E",X"61",X"6B",X"65",X"00",X"00",
		X"00",X"0E",X"18",X"39",X"FB",X"EE",X"19",X"41",
		X"00",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"00",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"FC",X"02",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"13",X"0C",X"C3",X"30",X"0C",
		X"C3",X"2A",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"AB",
		X"2A",X"0C",X"C3",X"00",X"FD",X"04",X"68",X"18",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"F0",X"0F",X"C3",X"30",
		X"0C",X"C3",X"F0",X"0F",X"C3",X"30",X"0C",X"C3",
		X"3F",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"15",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"1C",X"04",X"6B",X"00",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"3F",X"00",X"C3",X"30",
		X"0C",X"C3",X"F0",X"0F",X"C0",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"2A",X"0C",X"C3",X"30",X"0C",X"AB",X"2A",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"FF",X"FB",X"BF",
		X"3F",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"AC",X"56",X"95",X"0A",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"F0",X"FF",X"C3",X"30",
		X"0C",X"C3",X"F0",X"FF",X"C3",X"30",X"0C",X"C3",
		X"FF",X"0F",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"15",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"1C",X"00",X"FD",X"04",X"68",X"18",
		X"AC",X"56",X"60",X"59",X"30",X"0C",X"C3",X"70",
		X"55",X"FD",X"55",X"F5",X"57",X"D5",X"5F",X"55",
		X"7F",X"55",X"FD",X"55",X"05",X"C3",X"30",X"0C",
		X"C3",X"F0",X"0B",X"C0",X"30",X"0C",X"C3",X"2F",
		X"00",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"2A",X"0C",X"C3",
		X"B0",X"AA",X"AA",X"2A",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"BF",X"91",X"F4",X"46",X"D2",X"0B",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"AC",X"C2",X"B0",
		X"AA",X"AA",X"AA",X"AA",X"C2",X"B0",X"0A",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"AC",X"FE",X"FF",X"3F",X"C0",X"30",
		X"AC",X"FE",X"FF",X"3F",X"C0",X"B0",X"FA",X"FF",
		X"FF",X"00",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"57",X"55",X"05",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"96",X"15",
		X"58",X"6B",X"B0",X"AE",X"30",X"0C",X"C3",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"0F",X"C3",X"30",X"0C",
		X"C3",X"30",X"FC",X"03",X"30",X"0C",X"FF",X"00",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"FC",X"BF",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"00",X"FD",X"04",X"68",X"18",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"F0",
		X"FF",X"AB",X"FF",X"0F",X"C3",X"6A",X"A5",X"56",
		X"2A",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"FC",X"4A",X"30",
		X"FC",X"C2",X"70",X"F4",X"C2",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"F0",X"AF",X"FE",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"BF",X"FA",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"F0",X"FF",
		X"FF",X"30",X"0C",X"C3",X"F0",X"FF",X"FF",X"30",
		X"0C",X"C3",X"FF",X"FF",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"15",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"EB",X"1A",X"AC",X"56",X"B0",
		X"A6",X"30",X"0C",X"C3",X"70",X"55",X"FD",X"55",
		X"F5",X"57",X"D5",X"5F",X"55",X"7F",X"55",X"FD",
		X"55",X"05",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"BF",X"00",X"FC",X"02",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"6C",X"FC",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"F0",
		X"AF",X"FE",X"EA",X"0F",X"AB",X"AA",X"AA",X"AA",
		X"2A",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"F0",X"1B",X"BD",X"30",
		X"FC",X"C2",X"F0",X"2B",X"BD",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"00",X"FD",X"04",X"68",X"18",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"F0",X"AF",
		X"AB",X"95",X"5A",X"55",X"6A",X"A5",X"56",X"AA",
		X"FE",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"FF",X"AF",X"FE",X"30",X"0C",
		X"C3",X"FF",X"AF",X"FE",X"30",X"0C",X"FF",X"BF",
		X"FA",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"AB",X"95",
		X"0A",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"E9",X"1A",X"58",X"41",X"B0",X"AE",X"30",X"0C",
		X"C3",X"B0",X"AE",X"FE",X"AA",X"FE",X"AB",X"EA",
		X"AF",X"AB",X"BF",X"AA",X"FF",X"AA",X"0E",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"7F",X"05",
		X"C0",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"BC",X"BC",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"B0",X"FA",X"AB",X"BF",
		X"0A",X"AB",X"95",X"5A",X"A9",X"2A",X"0C",X"C3",
		X"12",X"5C",X"C2",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"BF",X"04",X"C3",X"2F",X"FC",X"C2",X"2F",
		X"0C",X"47",X"3F",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"B0",X"AA",
		X"AA",X"95",X"5A",X"A9",X"6A",X"A5",X"56",X"AA",
		X"AA",X"C2",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"0F",X"3F",X"AC",X"FE",X"30",X"0C",
		X"0F",X"3F",X"AC",X"FE",X"30",X"3C",X"FC",X"B0",
		X"FA",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"00",X"FD",X"04",X"68",X"18",
		X"C3",X"30",X"0C",X"C3",X"15",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"EB",X"1A",X"04",
		X"69",X"B0",X"A6",X"30",X"0C",X"C3",X"70",X"55",
		X"FD",X"55",X"F5",X"57",X"D5",X"5F",X"55",X"7F",
		X"55",X"FD",X"55",X"05",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"50",X"FD",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"6C",X"FC",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"70",X"A5",X"FE",X"EA",X"0F",X"AB",X"6A",
		X"A5",X"56",X"2A",X"0C",X"4B",X"92",X"54",X"96",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"6F",X"04",
		X"C3",X"F0",X"0B",X"BF",X"30",X"0C",X"4B",X"2F",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"AA",X"65",X"A9",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"65",X"A9",X"FF",
		X"FF",X"FF",X"FF",X"0F",X"C3",X"30",X"0C",X"C3",
		X"30",X"AC",X"FE",X"30",X"0C",X"C3",X"30",X"AC",
		X"FE",X"30",X"0C",X"C3",X"B0",X"FA",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"15",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"E9",X"1A",X"A4",
		X"41",X"B0",X"AE",X"30",X"0C",X"C3",X"B0",X"AA",
		X"FF",X"BA",X"FA",X"AB",X"FA",X"AF",X"AA",X"BF",
		X"AE",X"FE",X"BA",X"0A",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"C0",X"6B",X"01",X"2F",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"BC",X"BC",X"30",
		X"0C",X"C3",X"30",X"00",X"FD",X"04",X"68",X"18",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"B0",X"5A",
		X"A9",X"BF",X"0A",X"AB",X"95",X"5A",X"A9",X"2A",
		X"0C",X"4B",X"A3",X"94",X"97",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"FF",X"FB",X"BE",X"2F",X"FC",
		X"C3",X"EF",X"FB",X"BE",X"3F",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"AC",X"69",X"9A",X"A6",X"69",
		X"96",X"AA",X"1A",X"96",X"65",X"59",X"96",X"65",
		X"59",X"86",X"AA",X"5A",X"9A",X"A6",X"69",X"9A",
		X"06",X"C3",X"30",X"0C",X"C3",X"30",X"AC",X"FE",
		X"30",X"0C",X"C3",X"30",X"AC",X"FE",X"30",X"0C",
		X"C3",X"B0",X"FA",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"AC",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"15",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"EB",X"1A",X"04",X"69",X"B0",X"A6",
		X"30",X"0C",X"C3",X"70",X"55",X"FD",X"55",X"F5",
		X"57",X"D5",X"5F",X"55",X"7F",X"55",X"FD",X"55",
		X"05",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"03",
		X"7F",X"10",X"04",X"C0",X"0F",X"C3",X"30",X"0C",
		X"C3",X"30",X"6C",X"FC",X"41",X"10",X"04",X"41",
		X"10",X"04",X"41",X"10",X"04",X"41",X"10",X"04",
		X"41",X"10",X"04",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"70",X"A5",
		X"FE",X"EA",X"0F",X"AB",X"6A",X"A5",X"56",X"2A",
		X"1C",X"58",X"81",X"15",X"58",X"11",X"0C",X"C3",
		X"30",X"0C",X"C3",X"00",X"FD",X"04",X"68",X"18",
		X"AF",X"04",X"C3",X"F0",X"0F",X"FF",X"30",X"0C",
		X"47",X"2F",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"5C",X"55",X"55",X"55",X"55",X"D6",X"FA",X"5A",
		X"69",X"9A",X"A6",X"69",X"9A",X"A6",X"D6",X"BB",
		X"5A",X"55",X"55",X"55",X"55",X"05",X"C3",X"30",
		X"0C",X"C3",X"30",X"AC",X"FE",X"30",X"0C",X"C3",
		X"30",X"AC",X"FE",X"30",X"0C",X"C3",X"B0",X"FA",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"AB",X"AA",X"AA",X"AA",
		X"AA",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"E9",
		X"1A",X"A4",X"41",X"B0",X"AE",X"30",X"0C",X"C3",
		X"B0",X"AA",X"FF",X"AA",X"FE",X"AB",X"EA",X"AF",
		X"EA",X"BF",X"AA",X"FF",X"AA",X"0E",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"BC",X"81",X"65",X"05",
		X"20",X"F0",X"C2",X"30",X"0C",X"C3",X"30",X"BC",
		X"BC",X"FF",X"FB",X"BF",X"FF",X"FB",X"BF",X"FF",
		X"FB",X"BF",X"FF",X"FB",X"BF",X"FF",X"FB",X"07",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"B0",X"5A",X"A9",X"BF",X"0A",
		X"AB",X"95",X"5A",X"A9",X"2A",X"1C",X"04",X"41",
		X"10",X"44",X"11",X"0C",X"C3",X"30",X"0C",X"C3",
		X"7F",X"04",X"C3",X"EF",X"FF",X"FE",X"3F",X"0C",
		X"4B",X"3F",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"AC",X"AA",X"95",X"AA",X"56",X"D6",X"FA",X"5A",
		X"6A",X"A5",X"AA",X"6A",X"A5",X"AA",X"D6",X"BB",
		X"5A",X"95",X"AA",X"56",X"AA",X"0A",X"C3",X"30",
		X"0C",X"C3",X"30",X"AC",X"FE",X"30",X"0C",X"C3",
		X"30",X"AC",X"FE",X"30",X"0C",X"C3",X"B0",X"FA",
		X"C3",X"30",X"0C",X"00",X"FD",X"04",X"68",X"18",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"55",
		X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",
		X"EA",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0C",
		X"C3",X"30",X"0C",X"C3",X"EB",X"1A",X"04",X"69",
		X"B0",X"A6",X"30",X"0C",X"C3",X"70",X"55",X"FD",
		X"55",X"F5",X"57",X"D5",X"5F",X"55",X"7F",X"55",
		X"FD",X"55",X"05",X"C3",X"30",X"0C",X"C3",X"30",
		X"F0",X"83",X"81",X"65",X"05",X"20",X"08",X"FC",
		X"30",X"0C",X"C3",X"30",X"6C",X"FC",X"6F",X"60",
		X"04",X"46",X"60",X"04",X"46",X"60",X"04",X"C6",
		X"6F",X"2C",X"56",X"F0",X"06",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"70",X"A5",X"FE",X"EA",X"0F",X"AB",X"6A",X"A5",
		X"56",X"2A",X"1C",X"58",X"81",X"15",X"58",X"11",
		X"0C",X"C3",X"30",X"0C",X"C3",X"F0",X"0B",X"BF",
		X"3F",X"FC",X"C2",X"FF",X"0F",X"BF",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"AC",X"69",X"55",
		X"55",X"55",X"96",X"AA",X"5A",X"AA",X"6A",X"A9",
		X"96",X"AA",X"AA",X"96",X"AA",X"5A",X"55",X"55",
		X"55",X"9A",X"06",X"C3",X"30",X"0C",X"C3",X"30",
		X"AC",X"FE",X"30",X"0C",X"C3",X"30",X"AC",X"FE",
		X"30",X"0C",X"C3",X"B0",X"FA",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"00",X"00",X"00",
		X"00",X"00",X"55",X"55",X"55",X"55",X"A5",X"AA",
		X"AA",X"AA",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"30",X"0C",X"C3",X"E9",X"1A",X"A4",X"41",
		X"B0",X"AE",X"30",X"0C",X"C3",X"B0",X"AE",X"FE",
		X"BA",X"FA",X"AB",X"FA",X"AF",X"AA",X"BF",X"AE",
		X"FE",X"AA",X"0E",X"C3",X"30",X"0C",X"C3",X"C0",
		X"1B",X"04",X"41",X"00",X"FD",X"04",X"68",X"18",
		X"10",X"04",X"41",X"00",X"03",X"30",X"0C",X"C3",
		X"30",X"BC",X"BC",X"BF",X"F1",X"1A",X"8B",X"B1",
		X"18",X"8B",X"B1",X"18",X"C1",X"BB",X"58",X"46",
		X"F0",X"07",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"B0",X"5A",X"A9",
		X"BF",X"0A",X"AB",X"95",X"5A",X"A9",X"2A",X"1C",
		X"04",X"41",X"10",X"44",X"11",X"0C",X"C3",X"30",
		X"0C",X"C3",X"70",X"F4",X"FE",X"30",X"FC",X"C2",
		X"F0",X"FF",X"4B",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"AC",X"69",X"9A",X"AA",X"6A",X"16",
		X"A5",X"5A",X"AA",X"61",X"A9",X"56",X"65",X"A8",
		X"56",X"95",X"5A",X"9A",X"AA",X"6A",X"9A",X"06",
		X"C3",X"30",X"0C",X"C3",X"30",X"AC",X"FE",X"30",
		X"0C",X"C3",X"30",X"AC",X"FE",X"30",X"0C",X"C3",
		X"B0",X"FA",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"03",X"00",X"00",X"00",X"00",
		X"00",X"54",X"55",X"55",X"55",X"55",X"A5",X"AA",
		X"AA",X"FA",X"FF",X"FF",X"0F",X"C3",X"30",X"0C",
		X"C3",X"EB",X"1A",X"04",X"69",X"B0",X"A6",X"30",
		X"0C",X"C3",X"70",X"55",X"FD",X"55",X"F5",X"57",
		X"D5",X"5F",X"55",X"7F",X"55",X"FD",X"55",X"05",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"07",X"96",
		X"65",X"59",X"01",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"6C",X"FC",X"6F",X"60",X"2C",X"C6",X"62",
		X"2C",X"C6",X"62",X"2C",X"C6",X"6F",X"19",X"56",
		X"F0",X"06",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"0C",X"C3",X"70",X"A5",X"FE",
		X"EA",X"0F",X"AB",X"00",X"FD",X"04",X"68",X"18",
		X"6A",X"A5",X"56",X"2A",X"1C",X"58",X"81",X"15",
		X"58",X"11",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"FC",X"BF",X"30",X"FC",X"C2",X"F0",X"FB",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"5C",
		X"A9",X"69",X"55",X"55",X"29",X"55",X"55",X"55",
		X"55",X"51",X"54",X"55",X"55",X"14",X"90",X"52",
		X"55",X"55",X"55",X"6A",X"05",X"C3",X"30",X"0C",
		X"C3",X"30",X"AC",X"FE",X"30",X"0C",X"C3",X"30",
		X"AC",X"FE",X"30",X"0C",X"C3",X"B0",X"FA",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"55",X"55",X"55",X"55",X"55",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"E9",X"1A",
		X"A4",X"41",X"B0",X"AE",X"30",X"0C",X"C3",X"B0",
		X"4A",X"D3",X"34",X"4D",X"D3",X"34",X"4D",X"D3",
		X"34",X"4D",X"D3",X"B4",X"0A",X"C3",X"30",X"0C",
		X"C3",X"30",X"0C",X"07",X"96",X"45",X"58",X"01",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"BC",X"BC",
		X"BF",X"11",X"18",X"81",X"11",X"18",X"81",X"11",
		X"18",X"C1",X"1B",X"04",X"41",X"F0",X"07",X"30",
		X"0C",X"C3",X"30",X"0C",X"FC",X"30",X"0C",X"FF",
		X"3F",X"0C",X"C3",X"3F",X"F0",X"C3",X"30",X"0C",
		X"FF",X"C0",X"0F",X"C3",X"FF",X"0F",X"C3",X"30",
		X"0C",X"C3",X"B0",X"5A",X"A9",X"BF",X"0A",X"AB",
		X"95",X"5A",X"A9",X"2A",X"1C",X"04",X"41",X"10",
		X"44",X"11",X"0C",X"C3",X"30",X"0C",X"C3",X"F0",
		X"FF",X"4B",X"FF",X"FB",X"BF",X"BF",X"F4",X"FF",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"AC",
		X"AA",X"AA",X"5A",X"A9",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"6A",X"9A",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"6A",X"A5",X"69",X"9A",X"06",X"C3",X"30",X"0C",
		X"C3",X"30",X"AC",X"00",X"FD",X"04",X"68",X"18",
		X"FE",X"30",X"0C",X"C3",X"30",X"AC",X"FE",X"30",
		X"0C",X"C3",X"B0",X"FA",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"EB",X"1A",X"04",X"69",X"B0",
		X"A6",X"30",X"0C",X"C3",X"70",X"05",X"C3",X"FE",
		X"EF",X"FF",X"FE",X"EF",X"FF",X"FE",X"EF",X"C3",
		X"70",X"05",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"07",X"84",X"65",X"59",X"01",X"0C",X"C3",X"30",
		X"0C",X"C3",X"30",X"6C",X"FC",X"EF",X"FF",X"FE",
		X"EF",X"FF",X"FE",X"EF",X"FF",X"FE",X"EF",X"FF",
		X"FE",X"EF",X"FF",X"06",X"30",X"0C",X"C3",X"0C",
		X"F3",X"03",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"CC",X"FF",X"33",X"0C",X"C3",X"00",X"3F",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"0C",X"C3",X"70",
		X"A5",X"FE",X"EA",X"0F",X"AB",X"6A",X"A5",X"56",
		X"2A",X"1C",X"58",X"81",X"15",X"58",X"11",X"0C",
		X"C3",X"30",X"0C",X"C3",X"F0",X"0F",X"C3",X"52",
		X"24",X"05",X"12",X"0C",X"FF",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"5C",X"55",X"55",X"55",
		X"55",X"15",X"55",X"A9",X"95",X"AA",X"AA",X"AA",
		X"1A",X"54",X"41",X"55",X"55",X"55",X"55",X"05",
		X"95",X"0A",X"C3",X"30",X"CC",X"30",X"8C",X"FA",
		X"FF",X"3F",X"C3",X"30",X"8C",X"FA",X"FF",X"3F",
		X"C3",X"30",X"EA",X"FF",X"FF",X"0C",X"C3",X"C0",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"C3",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"15",X"0C",X"C3",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"E9",X"1A",X"A4",X"41",X"B0",
		X"AE",X"30",X"0C",X"C3",X"70",X"F5",X"FB",X"BF",
		X"AF",X"AA",X"AA",X"00",X"FD",X"04",X"68",X"18",
		X"AA",X"AA",X"AA",X"FA",X"FB",X"7F",X"05",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"07",X"84",X"65",
		X"59",X"01",X"0C",X"C3",X"30",X"0C",X"C3",X"30",
		X"BC",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"07",X"30",X"0C",X"33",X"08",X"82",X"20",X"08",
		X"82",X"20",X"08",X"82",X"20",X"08",X"82",X"20",
		X"08",X"82",X"20",X"08",X"82",X"20",X"08",X"82",
		X"20",X"08",X"03",X"C3",X"B0",X"5A",X"A9",X"BF",
		X"0A",X"AB",X"AA",X"AA",X"AA",X"2A",X"1C",X"04",
		X"41",X"10",X"44",X"11",X"0C",X"C3",X"30",X"0C",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"0F",X"C3",X"30",X"0C",X"C3",
		X"30",X"5C",X"14",X"45",X"51",X"14",X"45",X"51",
		X"14",X"45",X"51",X"14",X"45",X"51",X"14",X"45",
		X"51",X"14",X"45",X"51",X"14",X"45",X"01",X"C3",
		X"30",X"83",X"20",X"08",X"82",X"20",X"08",X"82",
		X"20",X"08",X"82",X"20",X"08",X"82",X"20",X"08",
		X"82",X"20",X"08",X"82",X"30",X"30",X"0C",X"C3",
		X"30",X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",
		X"03",X"00",X"00",X"00",X"00",X"00",X"C3",X"15",
		X"0C",X"C3",X"30",X"0C",X"C3",X"30",X"0C",X"C3",
		X"EB",X"1A",X"04",X"7A",X"69",X"70",X"70",X"65",
		X"64",X"52",X"61",X"77",X"18",X"40",X"FB",X"EE",
		X"19",X"02",X"00",X"F7",X"1A",X"21",X"E6",X"20",
		X"35",X"53",X"0B",X"21",X"0E",X"F3",X"17",X"90",
		X"05",X"CD",X"57",X"E6",X"52",X"35",X"53",X"1B",
		X"E3",X"32",X"2B",X"30",X"11",X"00",X"07",X"90",
		X"20",X"2B",X"30",X"11",X"00",X"08",X"2B",X"32",
		X"21",X"30",X"E9",X"E9",X"99",X"30",X"99",X"32",
		X"2B",X"32",X"21",X"34",X"5E",X"24",X"21",X"36",
		X"5E",X"25",X"21",X"00",X"FD",X"04",X"68",X"18",
		X"38",X"2B",X"28",X"11",X"E1",X"04",X"2B",X"22",
		X"59",X"FB",X"2B",X"30",X"21",X"32",X"7F",X"00",
		X"93",X"32",X"5E",X"26",X"B4",X"CB",X"93",X"28",
		X"93",X"30",X"21",X"30",X"35",X"72",X"41",X"21",
		X"38",X"FF",X"2B",X"3A",X"CD",X"F0",X"1A",X"0E",
		X"B8",X"3C",X"82",X"FF",X"5E",X"2B",X"99",X"3E",
		X"35",X"53",X"6B",X"11",X"FF",X"7F",X"2B",X"3E",
		X"1A",X"0E",X"2B",X"3C",X"1A",X"41",X"35",X"56",
		X"8A",X"2B",X"30",X"21",X"42",X"B8",X"44",X"2B",
		X"42",X"21",X"46",X"99",X"48",X"2B",X"46",X"21",
		X"30",X"E6",X"01",X"90",X"73",X"59",X"00",X"2B",
		X"4A",X"1A",X"11",X"82",X"01",X"35",X"72",X"A0",
		X"11",X"00",X"02",X"99",X"42",X"2B",X"42",X"59",
		X"01",X"2B",X"4A",X"1A",X"11",X"82",X"02",X"35",
		X"72",X"B3",X"11",X"00",X"FE",X"99",X"42",X"2B",
		X"42",X"11",X"FF",X"FF",X"2B",X"4A",X"1A",X"11",
		X"82",X"80",X"35",X"72",X"CF",X"21",X"40",X"E3",
		X"10",X"2B",X"40",X"11",X"FF",X"05",X"B8",X"40",
		X"35",X"53",X"CD",X"11",X"FF",X"05",X"2B",X"40",
		X"90",X"DD",X"11",X"F8",X"FE",X"99",X"40",X"35",
		X"50",X"DD",X"21",X"40",X"E6",X"08",X"2B",X"40",
		X"1A",X"11",X"82",X"40",X"35",X"72",X"EF",X"21",
		X"40",X"E6",X"40",X"35",X"53",X"ED",X"59",X"00",
		X"2B",X"40",X"FF",X"2B",X"4C",X"93",X"1B",X"FF",
		X"03",X"00",X"E1",X"CD",X"09",X"47",X"69",X"67",
		X"61",X"74",X"72",X"6F",X"6E",X"00",X"2B",X"4E",
		X"CD",X"1D",X"1A",X"0E",X"99",X"50",X"82",X"FF",
		X"2B",X"52",X"1A",X"0E",X"B8",X"52",X"35",X"72",
		X"15",X"FF",X"2B",X"54",X"CD",X"A1",X"21",X"56",
		X"AD",X"82",X"FE",X"5E",X"59",X"88",X"01",X"5E",
		X"5B",X"93",X"56",X"59",X"00",X"5E",X"58",X"5E",
		X"5A",X"21",X"58",X"00",X"FD",X"04",X"68",X"18",
		X"AD",X"2B",X"30",X"21",X"5A",X"AD",X"B8",X"30",
		X"2B",X"30",X"21",X"58",X"AD",X"5E",X"58",X"5E",
		X"5A",X"59",X"15",X"F0",X"58",X"F0",X"5A",X"93",
		X"58",X"93",X"5A",X"21",X"30",X"E6",X"01",X"2B",
		X"30",X"35",X"4D",X"47",X"21",X"5C",X"2B",X"5E",
		X"59",X"00",X"5E",X"58",X"21",X"56",X"AD",X"99",
		X"60",X"2B",X"60",X"21",X"5E",X"AD",X"99",X"60",
		X"F0",X"58",X"5E",X"58",X"5E",X"5A",X"93",X"5E",
		X"21",X"58",X"AD",X"8C",X"15",X"99",X"62",X"2B",
		X"62",X"21",X"5E",X"AD",X"F0",X"58",X"93",X"58",
		X"F0",X"5A",X"93",X"5A",X"93",X"5E",X"21",X"5E",
		X"AD",X"35",X"72",X"76",X"59",X"00",X"5E",X"5A",
		X"1A",X"58",X"F0",X"5A",X"21",X"56",X"E3",X"03",
		X"2B",X"56",X"FF",X"2B",X"64",X"CD",X"DA",X"11",
		X"FD",X"01",X"2B",X"58",X"21",X"40",X"99",X"40",
		X"1A",X"19",X"F0",X"58",X"93",X"59",X"F0",X"58",
		X"93",X"59",X"F0",X"58",X"93",X"59",X"F0",X"58",
		X"11",X"FC",X"01",X"2B",X"58",X"21",X"40",X"82",
		X"7F",X"F0",X"58",X"93",X"59",X"F0",X"58",X"93",
		X"59",X"F0",X"58",X"93",X"59",X"F0",X"58",X"59",
		X"0A",X"5E",X"2C",X"FF",X"2B",X"66",X"93",X"1B",
		X"FF",X"04",X"00",X"EF",X"CD",X"3E",X"75",X"11",
		X"80",X"20",X"2B",X"38",X"11",X"03",X"0B",X"2B",
		X"22",X"59",X"00",X"2B",X"68",X"21",X"68",X"E3",
		X"01",X"2B",X"68",X"59",X"3F",X"2B",X"6A",X"59",
		X"0C",X"2B",X"6C",X"CF",X"6E",X"93",X"39",X"59",
		X"03",X"2B",X"6A",X"59",X"08",X"2B",X"6C",X"CF",
		X"6E",X"93",X"39",X"21",X"38",X"35",X"53",X"0F",
		X"11",X"00",X"74",X"F0",X"18",X"93",X"19",X"35",
		X"4D",X"35",X"63",X"FF",X"2B",X"70",X"CD",X"86",
		X"21",X"68",X"E9",X"5E",X"24",X"21",X"38",X"B8",
		X"68",X"2B",X"58",X"00",X"FD",X"04",X"68",X"18",
		X"2B",X"26",X"59",X"15",X"5E",X"25",X"B4",X"F3",
		X"59",X"80",X"B8",X"68",X"E9",X"5E",X"24",X"21",
		X"38",X"99",X"68",X"2B",X"5A",X"2B",X"26",X"21",
		X"6C",X"5E",X"25",X"B4",X"F3",X"21",X"68",X"E6",
		X"08",X"35",X"56",X"85",X"2B",X"52",X"21",X"5A",
		X"E6",X"01",X"2B",X"5A",X"21",X"6A",X"F0",X"58",
		X"F0",X"5A",X"93",X"58",X"21",X"52",X"90",X"6C",
		X"FF",X"2B",X"6E",X"CD",X"E8",X"75",X"11",X"0F",
		X"0E",X"2B",X"72",X"CF",X"74",X"21",X"76",X"FC",
		X"78",X"35",X"3F",X"A1",X"21",X"78",X"2B",X"76",
		X"CF",X"3A",X"90",X"A3",X"21",X"38",X"E3",X"0C",
		X"2B",X"38",X"11",X"58",X"02",X"2B",X"72",X"CF",
		X"74",X"21",X"7A",X"FC",X"78",X"35",X"3F",X"BD",
		X"21",X"78",X"2B",X"7A",X"CF",X"3A",X"90",X"BF",
		X"21",X"38",X"E3",X"06",X"2B",X"38",X"59",X"3C",
		X"2B",X"72",X"CF",X"74",X"21",X"7C",X"FC",X"78",
		X"35",X"3F",X"D8",X"21",X"78",X"2B",X"7C",X"CF",
		X"3A",X"90",X"DA",X"21",X"38",X"E3",X"0C",X"2B",
		X"38",X"59",X"06",X"2B",X"72",X"CF",X"74",X"CF",
		X"3A",X"63",X"FF",X"2B",X"7E",X"93",X"1B",X"FF",
		X"05",X"00",X"E6",X"CD",X"17",X"59",X"30",X"2B",
		X"78",X"21",X"81",X"B8",X"72",X"35",X"50",X"14",
		X"2B",X"81",X"93",X"78",X"B8",X"72",X"35",X"53",
		X"0B",X"21",X"78",X"FF",X"2B",X"74",X"CD",X"32",
		X"75",X"2B",X"83",X"21",X"83",X"AD",X"2B",X"78",
		X"35",X"3F",X"30",X"93",X"83",X"CF",X"3A",X"E3",
		X"06",X"2B",X"38",X"90",X"1E",X"63",X"FF",X"2B",
		X"85",X"CD",X"DF",X"11",X"D0",X"74",X"2B",X"58",
		X"59",X"00",X"2B",X"60",X"21",X"87",X"2B",X"89",
		X"21",X"8B",X"B8",X"8D",X"2B",X"52",X"99",X"52",
		X"2B",X"52",X"11",X"00",X"0A",X"99",X"52",X"7F",
		X"35",X"2B",X"52",X"00",X"FD",X"04",X"68",X"18",
		X"59",X"C5",X"99",X"52",X"2B",X"30",X"1A",X"61",
		X"F0",X"58",X"93",X"58",X"21",X"89",X"99",X"8F",
		X"2B",X"89",X"99",X"60",X"2B",X"60",X"93",X"30",
		X"21",X"30",X"35",X"72",X"5C",X"1A",X"61",X"F0",
		X"58",X"93",X"58",X"21",X"89",X"99",X"91",X"2B",
		X"89",X"99",X"60",X"2B",X"60",X"1A",X"58",X"35",
		X"72",X"73",X"11",X"ED",X"01",X"2B",X"24",X"11",
		X"D1",X"74",X"2B",X"26",X"E6",X"01",X"AD",X"2B",
		X"28",X"1A",X"47",X"2B",X"52",X"11",X"D5",X"74",
		X"AD",X"E3",X"30",X"B8",X"52",X"2B",X"52",X"11",
		X"D4",X"74",X"AD",X"2B",X"87",X"11",X"EC",X"74",
		X"AD",X"B8",X"87",X"82",X"FF",X"8C",X"80",X"E6",
		X"80",X"2B",X"87",X"11",X"11",X"01",X"2B",X"5E",
		X"1A",X"09",X"82",X"01",X"35",X"3F",X"BE",X"1A",
		X"47",X"F0",X"5E",X"11",X"38",X"40",X"2B",X"22",
		X"B4",X"FA",X"21",X"24",X"2B",X"5E",X"21",X"28",
		X"2B",X"60",X"21",X"52",X"B8",X"60",X"F0",X"5E",
		X"FF",X"2B",X"93",X"93",X"1B",X"FF",X"06",X"00",
		X"DF",X"CD",X"A7",X"75",X"59",X"00",X"2B",X"62",
		X"2B",X"76",X"2B",X"7A",X"2B",X"7C",X"CF",X"95",
		X"21",X"8D",X"35",X"53",X"2E",X"21",X"3E",X"B8",
		X"97",X"35",X"53",X"1D",X"21",X"3E",X"2B",X"97",
		X"59",X"0F",X"CF",X"99",X"59",X"00",X"2B",X"3E",
		X"2B",X"9B",X"11",X"00",X"74",X"2B",X"8D",X"2B",
		X"8B",X"B8",X"8B",X"35",X"56",X"73",X"21",X"9B",
		X"99",X"8B",X"8C",X"6D",X"2B",X"9B",X"82",X"1F",
		X"E3",X"28",X"99",X"8B",X"2B",X"8B",X"1A",X"9C",
		X"82",X"03",X"E3",X"01",X"2B",X"30",X"99",X"30",
		X"99",X"30",X"E9",X"2B",X"30",X"21",X"91",X"2B",
		X"8F",X"35",X"53",X"5D",X"99",X"30",X"90",X"71",
		X"35",X"56",X"64",X"B8",X"30",X"90",X"71",X"21",
		X"9B",X"35",X"50",X"00",X"FD",X"04",X"68",X"18",
		X"6D",X"21",X"30",X"90",X"71",X"59",X"00",X"B8",
		X"30",X"2B",X"91",X"CF",X"93",X"21",X"8F",X"E9",
		X"E9",X"E9",X"2B",X"48",X"E9",X"2B",X"44",X"CF",
		X"4C",X"CF",X"66",X"CF",X"9D",X"CF",X"9F",X"11",
		X"B5",X"B9",X"99",X"3E",X"35",X"56",X"91",X"2B",
		X"62",X"21",X"3E",X"2B",X"81",X"11",X"01",X"08",
		X"2B",X"38",X"59",X"3F",X"2B",X"36",X"CF",X"7E",
		X"21",X"62",X"35",X"3F",X"0B",X"63",X"FF",X"2B",
		X"A1",X"CD",X"B7",X"02",X"40",X"40",X"40",X"28",
		X"3C",X"3C",X"28",X"40",X"40",X"40",X"00",X"2B",
		X"A3",X"CD",X"C5",X"03",X"28",X"14",X"14",X"3F",
		X"3F",X"14",X"14",X"28",X"00",X"2B",X"A5",X"CD",
		X"D5",X"02",X"28",X"14",X"14",X"14",X"28",X"28",
		X"14",X"14",X"14",X"28",X"00",X"2B",X"A7",X"11",
		X"A0",X"08",X"2B",X"1A",X"FF",X"08",X"A0",X"52",
		X"CD",X"B0",X"00",X"40",X"40",X"40",X"40",X"28",
		X"14",X"14",X"14",X"14",X"28",X"40",X"40",X"40",
		X"40",X"00",X"2B",X"A9",X"CD",X"C4",X"00",X"40",
		X"40",X"40",X"40",X"15",X"15",X"15",X"15",X"15",
		X"15",X"40",X"40",X"40",X"40",X"00",X"2B",X"AB",
		X"CD",X"EB",X"11",X"2E",X"01",X"2B",X"24",X"59",
		X"20",X"5E",X"26",X"11",X"00",X"0A",X"2B",X"5A",
		X"11",X"51",X"40",X"2B",X"22",X"21",X"5A",X"7F",
		X"08",X"99",X"8D",X"5E",X"27",X"B4",X"FA",X"93",
		X"5A",X"35",X"72",X"DB",X"FF",X"2B",X"9F",X"93",
		X"1B",X"FF",X"09",X"A0",X"38",X"CD",X"B8",X"11",
		X"F7",X"0B",X"2B",X"AD",X"11",X"6B",X"0C",X"2B",
		X"AF",X"59",X"00",X"F0",X"AF",X"93",X"AF",X"1A",
		X"AF",X"8C",X"76",X"35",X"72",X"AA",X"FF",X"2B",
		X"B1",X"CD",X"D1",X"59",X"00",X"F0",X"AF",X"1A",
		X"8E",X"99",X"AD",X"2B",X"AF",X"59",X"3C",X"F0",
		X"AF",X"1A",X"41",X"00",X"FD",X"04",X"68",X"18",
		X"99",X"8D",X"2B",X"8D",X"FF",X"2B",X"95",X"93",
		X"1B",X"FF",X"0A",X"A0",X"41",X"CD",X"DA",X"75",
		X"11",X"D9",X"01",X"AD",X"8C",X"FF",X"2B",X"60",
		X"1A",X"43",X"99",X"60",X"2B",X"60",X"11",X"D8",
		X"01",X"2B",X"56",X"21",X"A3",X"2B",X"5C",X"CF",
		X"64",X"21",X"A5",X"2B",X"5C",X"CF",X"64",X"21",
		X"60",X"B8",X"4A",X"2B",X"60",X"21",X"A7",X"2B",
		X"5C",X"CF",X"64",X"21",X"A9",X"2B",X"5C",X"CF",
		X"64",X"21",X"AB",X"2B",X"5C",X"CF",X"64",X"63",
		X"FF",X"2B",X"9D",X"93",X"1B",X"FF",X"0B",X"A0",
		X"4C",X"CD",X"E5",X"75",X"59",X"30",X"2B",X"34",
		X"21",X"34",X"5E",X"24",X"5E",X"25",X"11",X"00",
		X"08",X"2B",X"28",X"11",X"E1",X"04",X"2B",X"22",
		X"B4",X"CB",X"93",X"28",X"1A",X"28",X"8C",X"A0",
		X"35",X"72",X"B5",X"59",X"3F",X"2B",X"36",X"11",
		X"07",X"08",X"2B",X"38",X"59",X"3A",X"CF",X"3A",
		X"E3",X"12",X"2B",X"38",X"59",X"2E",X"CF",X"3A",
		X"E3",X"1F",X"2B",X"38",X"21",X"4E",X"CF",X"85",
		X"59",X"3C",X"2B",X"50",X"CF",X"54",X"63",X"FF",
		X"2B",X"B3",X"93",X"1B",X"FF",X"0C",X"A0",X"59",
		X"CD",X"F2",X"2B",X"36",X"21",X"97",X"2B",X"81",
		X"E3",X"01",X"35",X"53",X"AC",X"FF",X"75",X"11",
		X"7C",X"08",X"2B",X"38",X"11",X"0F",X"0E",X"2B",
		X"72",X"CF",X"74",X"CF",X"3A",X"E3",X"06",X"2B",
		X"38",X"59",X"3A",X"CF",X"3A",X"E3",X"06",X"2B",
		X"38",X"11",X"58",X"02",X"2B",X"72",X"CF",X"74",
		X"CF",X"3A",X"E3",X"06",X"2B",X"38",X"59",X"3C",
		X"2B",X"72",X"CF",X"74",X"CF",X"3A",X"E3",X"06",
		X"2B",X"38",X"59",X"2E",X"CF",X"3A",X"E3",X"06",
		X"2B",X"38",X"59",X"06",X"2B",X"72",X"CF",X"74",
		X"CF",X"3A",X"63",X"FF",X"2B",X"99",X"93",X"1B",
		X"FF",X"0D",X"A0",X"00",X"FD",X"04",X"68",X"18",
		X"56",X"CD",X"EF",X"75",X"11",X"35",X"14",X"2B",
		X"38",X"CD",X"B2",X"47",X"41",X"4D",X"45",X"20",
		X"4F",X"56",X"45",X"52",X"00",X"CF",X"85",X"11",
		X"11",X"01",X"2B",X"5E",X"E3",X"20",X"2B",X"B5",
		X"59",X"01",X"2B",X"50",X"21",X"5E",X"AD",X"82",
		X"80",X"35",X"72",X"CD",X"59",X"01",X"90",X"D0",
		X"11",X"FF",X"FF",X"2B",X"30",X"CF",X"54",X"21",
		X"B5",X"AD",X"B8",X"30",X"F0",X"B5",X"21",X"5E",
		X"AD",X"99",X"30",X"F0",X"5E",X"82",X"FF",X"35",
		X"72",X"D2",X"59",X"1E",X"2B",X"50",X"CF",X"54",
		X"63",X"FF",X"2B",X"B7",X"93",X"1B",X"FF",X"0E",
		X"A0",X"5B",X"CD",X"F4",X"75",X"11",X"77",X"40",
		X"2B",X"58",X"11",X"00",X"10",X"2B",X"5A",X"CD",
		X"BF",X"1A",X"58",X"8C",X"FA",X"35",X"3F",X"B8",
		X"59",X"01",X"90",X"BA",X"59",X"06",X"99",X"58",
		X"2B",X"58",X"FF",X"2B",X"52",X"21",X"58",X"7F",
		X"00",X"5E",X"24",X"CF",X"52",X"7F",X"00",X"5E",
		X"25",X"CF",X"52",X"7F",X"00",X"5E",X"26",X"CF",
		X"52",X"11",X"C0",X"06",X"2B",X"22",X"B4",X"F2",
		X"21",X"5A",X"2B",X"28",X"E3",X"04",X"2B",X"5A",
		X"11",X"D4",X"04",X"2B",X"22",X"B4",X"FF",X"1A",
		X"5B",X"8C",X"20",X"35",X"72",X"C1",X"63",X"FF",
		X"2B",X"B9",X"93",X"1B",X"FF",X"0F",X"A0",X"54",
		X"CF",X"B3",X"11",X"00",X"74",X"2B",X"8D",X"2B",
		X"8B",X"11",X"FF",X"7F",X"2B",X"97",X"59",X"00",
		X"2B",X"3E",X"2B",X"81",X"2B",X"46",X"2B",X"44",
		X"2B",X"40",X"2B",X"9B",X"2B",X"87",X"2B",X"8F",
		X"2B",X"91",X"CF",X"93",X"CF",X"9F",X"CF",X"B9",
		X"11",X"35",X"14",X"2B",X"38",X"CD",X"D7",X"47",
		X"45",X"54",X"20",X"52",X"45",X"41",X"44",X"59",
		X"00",X"CF",X"85",X"CF",X"70",X"CF",X"B9",X"CF",
		X"B1",X"11",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"79",X"2B",X"42",X"1A",X"0E",X"2B",X"3C",X"CF",
		X"A1",X"CF",X"B7",X"59",X"3F",X"CF",X"99",X"90",
		X"A0",X"00",X"52",X"61",X"63",X"65",X"72",X"00",
		X"00",X"00",X"C1",X"18",X"4C",X"FB",X"EE",X"19",
		X"02",X"00",X"EF",X"CD",X"E8",X"75",X"59",X"00",
		X"2B",X"30",X"2B",X"32",X"B8",X"34",X"35",X"56",
		X"12",X"2B",X"34",X"59",X"01",X"2B",X"30",X"59",
		X"00",X"B8",X"36",X"35",X"56",X"21",X"2B",X"36",
		X"21",X"30",X"8C",X"01",X"2B",X"30",X"59",X"07",
		X"2B",X"38",X"11",X"00",X"06",X"2B",X"22",X"11",
		X"00",X"02",X"2B",X"3A",X"11",X"00",X"C0",X"99",
		X"32",X"35",X"53",X"3E",X"21",X"32",X"E9",X"2B",
		X"32",X"90",X"4A",X"21",X"36",X"B4",X"F6",X"2B",
		X"36",X"21",X"38",X"E6",X"01",X"2B",X"38",X"21",
		X"34",X"B8",X"3A",X"35",X"50",X"59",X"2B",X"34",
		X"21",X"32",X"99",X"36",X"2B",X"32",X"21",X"3A",
		X"B4",X"F6",X"35",X"72",X"2D",X"21",X"38",X"8C",
		X"07",X"35",X"72",X"72",X"11",X"B9",X"04",X"2B",
		X"22",X"21",X"32",X"B4",X"FF",X"90",X"D7",X"21",
		X"38",X"8C",X"06",X"35",X"72",X"84",X"11",X"87",
		X"06",X"2B",X"22",X"21",X"32",X"B4",X"F6",X"90",
		X"D7",X"21",X"38",X"8C",X"05",X"35",X"72",X"96",
		X"11",X"6D",X"06",X"2B",X"22",X"21",X"32",X"B4",
		X"F5",X"90",X"D7",X"21",X"38",X"8C",X"04",X"35",
		X"72",X"A8",X"11",X"52",X"06",X"2B",X"22",X"21",
		X"32",X"B4",X"F5",X"90",X"D7",X"21",X"38",X"8C",
		X"03",X"35",X"72",X"BA",X"11",X"36",X"06",X"2B",
		X"22",X"21",X"32",X"B4",X"F4",X"90",X"D7",X"21",
		X"38",X"8C",X"02",X"35",X"72",X"CC",X"11",X"19",
		X"06",X"2B",X"22",X"21",X"32",X"B4",X"F4",X"90",
		X"D7",X"21",X"38",X"8C",X"01",X"35",X"72",X"D7",
		X"21",X"32",X"B4",X"00",X"FD",X"04",X"68",X"18",
		X"F6",X"2B",X"32",X"21",X"30",X"35",X"3F",X"E4",
		X"59",X"00",X"B8",X"32",X"90",X"E6",X"21",X"32",
		X"63",X"FF",X"2B",X"3C",X"93",X"1B",X"FF",X"03",
		X"00",X"EB",X"CD",X"E4",X"75",X"11",X"00",X"08",
		X"2B",X"3E",X"59",X"78",X"2B",X"40",X"59",X"A0",
		X"2B",X"42",X"2B",X"44",X"2B",X"46",X"59",X"00",
		X"2B",X"48",X"21",X"4A",X"2B",X"4C",X"59",X"3F",
		X"F0",X"3E",X"CF",X"4E",X"21",X"46",X"35",X"72",
		X"71",X"21",X"50",X"2B",X"34",X"2B",X"36",X"CF",
		X"3C",X"2B",X"52",X"21",X"54",X"E3",X"80",X"2B",
		X"34",X"2B",X"36",X"CF",X"3C",X"99",X"52",X"E6",
		X"08",X"35",X"53",X"44",X"59",X"00",X"90",X"6F",
		X"21",X"54",X"E6",X"20",X"2B",X"34",X"2B",X"36",
		X"CF",X"3C",X"99",X"52",X"2B",X"34",X"99",X"54",
		X"E6",X"20",X"2B",X"36",X"CF",X"3C",X"2B",X"56",
		X"99",X"56",X"2B",X"56",X"99",X"56",X"2B",X"56",
		X"B8",X"52",X"35",X"53",X"6D",X"59",X"00",X"90",
		X"6F",X"CF",X"58",X"90",X"73",X"CF",X"58",X"2B",
		X"46",X"F0",X"3E",X"21",X"44",X"E6",X"01",X"35",
		X"4D",X"9F",X"21",X"48",X"2B",X"56",X"21",X"4C",
		X"2B",X"48",X"59",X"00",X"B8",X"56",X"2B",X"4C",
		X"21",X"4C",X"35",X"3F",X"99",X"21",X"42",X"E6",
		X"01",X"2B",X"42",X"90",X"9F",X"21",X"40",X"E6",
		X"01",X"2B",X"40",X"2B",X"44",X"35",X"56",X"E0",
		X"21",X"54",X"99",X"4C",X"2B",X"54",X"21",X"50",
		X"99",X"48",X"2B",X"50",X"21",X"4C",X"35",X"53",
		X"BB",X"21",X"3E",X"E6",X"01",X"2B",X"3E",X"21",
		X"4C",X"35",X"56",X"C6",X"21",X"3E",X"E3",X"01",
		X"2B",X"3E",X"21",X"48",X"35",X"53",X"D2",X"11",
		X"00",X"FF",X"99",X"3E",X"2B",X"3E",X"21",X"48",
		X"35",X"56",X"DE",X"11",X"00",X"01",X"99",X"3E",
		X"2B",X"3E",X"90",X"00",X"FD",X"04",X"68",X"18",
		X"1A",X"CF",X"5A",X"63",X"FF",X"2B",X"5C",X"93",
		X"1B",X"FF",X"04",X"00",X"F0",X"CD",X"E4",X"75",
		X"11",X"00",X"08",X"2B",X"3E",X"59",X"78",X"2B",
		X"40",X"59",X"A0",X"2B",X"42",X"2B",X"44",X"59",
		X"01",X"2B",X"4C",X"59",X"00",X"2B",X"48",X"11",
		X"00",X"06",X"2B",X"22",X"59",X"00",X"2B",X"5E",
		X"59",X"20",X"2B",X"60",X"21",X"3E",X"AD",X"82",
		X"3F",X"B8",X"60",X"35",X"50",X"42",X"F0",X"3E",
		X"21",X"60",X"82",X"15",X"35",X"3F",X"3C",X"59",
		X"01",X"90",X"3E",X"59",X"02",X"99",X"5E",X"2B",
		X"5E",X"21",X"60",X"B4",X"F6",X"35",X"4D",X"23",
		X"F0",X"3E",X"21",X"5E",X"35",X"3F",X"83",X"1A",
		X"3F",X"82",X"01",X"2B",X"60",X"99",X"60",X"2B",
		X"60",X"21",X"3E",X"82",X"01",X"99",X"60",X"2B",
		X"60",X"CD",X"68",X"00",X"02",X"03",X"01",X"99",
		X"60",X"AD",X"99",X"5E",X"E6",X"01",X"2B",X"5E",
		X"21",X"5E",X"E6",X"03",X"35",X"50",X"83",X"2B",
		X"5E",X"21",X"3E",X"AD",X"E3",X"15",X"F0",X"3E",
		X"90",X"71",X"21",X"44",X"E6",X"01",X"35",X"4D",
		X"AB",X"21",X"48",X"2B",X"56",X"21",X"4C",X"2B",
		X"48",X"59",X"00",X"B8",X"56",X"2B",X"4C",X"21",
		X"4C",X"35",X"3F",X"A5",X"21",X"42",X"E6",X"01",
		X"2B",X"42",X"90",X"AB",X"21",X"40",X"E6",X"01",
		X"2B",X"40",X"2B",X"44",X"35",X"56",X"E2",X"21",
		X"4C",X"35",X"53",X"BB",X"21",X"3E",X"E6",X"01",
		X"2B",X"3E",X"21",X"4C",X"35",X"56",X"C6",X"21",
		X"3E",X"E3",X"01",X"2B",X"3E",X"21",X"48",X"35",
		X"53",X"D2",X"11",X"00",X"FF",X"99",X"3E",X"2B",
		X"3E",X"21",X"48",X"35",X"56",X"DE",X"11",X"00",
		X"01",X"99",X"3E",X"2B",X"3E",X"CF",X"4E",X"90",
		X"18",X"63",X"FF",X"2B",X"5A",X"11",X"1A",X"20",
		X"2B",X"62",X"93",X"00",X"FD",X"04",X"68",X"18",
		X"1B",X"FF",X"05",X"00",X"F6",X"CD",X"A4",X"1A",
		X"0E",X"B8",X"64",X"82",X"FF",X"2B",X"66",X"E6",
		X"3C",X"35",X"53",X"19",X"1A",X"11",X"82",X"80",
		X"35",X"3F",X"15",X"FF",X"59",X"0F",X"90",X"1B",
		X"59",X"3F",X"2B",X"68",X"75",X"21",X"6A",X"99",
		X"66",X"2B",X"6A",X"21",X"64",X"99",X"66",X"2B",
		X"64",X"11",X"F1",X"F1",X"99",X"6A",X"35",X"50",
		X"38",X"2B",X"6A",X"59",X"01",X"CF",X"6C",X"1A",
		X"63",X"FC",X"62",X"5E",X"63",X"1A",X"11",X"8C",
		X"77",X"35",X"72",X"4B",X"2B",X"6A",X"59",X"01",
		X"90",X"70",X"8C",X"0C",X"35",X"72",X"57",X"2B",
		X"6A",X"11",X"FF",X"FF",X"90",X"70",X"8C",X"06",
		X"35",X"72",X"63",X"2B",X"6A",X"11",X"C4",X"FF",
		X"90",X"70",X"8C",X"03",X"35",X"72",X"6E",X"2B",
		X"6A",X"59",X"3C",X"90",X"70",X"59",X"00",X"35",
		X"3F",X"7E",X"CF",X"6C",X"59",X"00",X"2B",X"6A",
		X"11",X"00",X"3A",X"2B",X"62",X"1A",X"11",X"88",
		X"0F",X"5E",X"11",X"11",X"5C",X"44",X"2B",X"6E",
		X"21",X"70",X"2B",X"72",X"11",X"58",X"02",X"CF",
		X"74",X"59",X"3C",X"CF",X"74",X"1A",X"63",X"CF",
		X"76",X"59",X"0A",X"CF",X"74",X"59",X"01",X"CF",
		X"74",X"63",X"FF",X"2B",X"4E",X"CD",X"EF",X"E6",
		X"20",X"2B",X"60",X"11",X"00",X"07",X"2B",X"78",
		X"21",X"60",X"E9",X"E9",X"99",X"60",X"99",X"78",
		X"2B",X"78",X"11",X"00",X"08",X"99",X"6E",X"2B",
		X"7A",X"59",X"00",X"5E",X"24",X"21",X"68",X"5E",
		X"25",X"21",X"6E",X"2B",X"28",X"E3",X"06",X"2B",
		X"6E",X"11",X"E1",X"04",X"2B",X"22",X"59",X"FB",
		X"2B",X"60",X"21",X"78",X"7F",X"00",X"93",X"78",
		X"5E",X"26",X"B4",X"CB",X"93",X"28",X"93",X"60",
		X"21",X"60",X"35",X"72",X"DB",X"FF",X"2B",X"76",
		X"93",X"1B",X"FF",X"00",X"FD",X"04",X"68",X"18",
		X"06",X"00",X"FE",X"CD",X"1D",X"75",X"2B",X"7C",
		X"59",X"30",X"2B",X"7E",X"21",X"72",X"B8",X"7C",
		X"35",X"50",X"17",X"2B",X"72",X"93",X"7E",X"B8",
		X"7C",X"35",X"53",X"0E",X"21",X"7E",X"CF",X"76",
		X"63",X"FF",X"2B",X"74",X"CD",X"3A",X"99",X"70",
		X"2B",X"70",X"35",X"53",X"2F",X"11",X"A0",X"05",
		X"99",X"70",X"2B",X"70",X"11",X"60",X"FA",X"99",
		X"70",X"35",X"50",X"39",X"2B",X"70",X"FF",X"2B",
		X"6C",X"CD",X"8E",X"75",X"59",X"00",X"2B",X"81",
		X"2B",X"83",X"2B",X"85",X"2B",X"52",X"2B",X"60",
		X"21",X"60",X"E3",X"01",X"2B",X"60",X"8C",X"40",
		X"35",X"3F",X"8C",X"21",X"81",X"2B",X"34",X"21",
		X"85",X"99",X"85",X"2B",X"36",X"CF",X"3C",X"99",
		X"50",X"2B",X"85",X"21",X"83",X"B8",X"52",X"99",
		X"54",X"2B",X"81",X"2B",X"34",X"2B",X"36",X"CF",
		X"3C",X"2B",X"83",X"21",X"85",X"2B",X"34",X"2B",
		X"36",X"CF",X"3C",X"2B",X"52",X"11",X"00",X"FE",
		X"99",X"83",X"99",X"52",X"35",X"56",X"4B",X"21",
		X"60",X"63",X"FF",X"2B",X"58",X"59",X"00",X"2B",
		X"6A",X"2B",X"70",X"2B",X"7E",X"1A",X"0E",X"2B",
		X"64",X"11",X"4C",X"FF",X"2B",X"50",X"11",X"C0",
		X"FE",X"2B",X"54",X"59",X"03",X"2B",X"4A",X"CF",
		X"5C",X"11",X"6C",X"FF",X"2B",X"50",X"11",X"9E",
		X"FF",X"2B",X"54",X"59",X"01",X"2B",X"4A",X"CF",
		X"5C",X"11",X"C4",X"FF",X"2B",X"50",X"11",X"00",
		X"FF",X"2B",X"54",X"59",X"01",X"2B",X"4A",X"CF",
		X"5C",X"11",X"C0",X"FE",X"2B",X"50",X"11",X"98",
		X"FE",X"2B",X"54",X"59",X"09",X"2B",X"4A",X"CF",
		X"5C",X"59",X"00",X"2B",X"50",X"11",X"9C",X"FF",
		X"2B",X"54",X"59",X"01",X"2B",X"4A",X"CF",X"5C",
		X"11",X"C4",X"FF",X"2B",X"50",X"59",X"00",X"2B",
		X"54",X"59",X"01",X"00",X"FD",X"04",X"68",X"18",
		X"2B",X"4A",X"CF",X"5C",X"90",X"9C",X"00",X"09",
		X"27",X"16",X"24",X"25",X"00",X"00",X"26",X"26",
		X"24",X"01",X"24",X"03",X"CB",X"F0",X"16",X"02",
		X"16",X"03",X"00",X"F3",X"25",X"26",X"48",X"24",
		X"41",X"00",X"00",X"4C",X"4C",X"00",X"00",X"3F",
		X"28",X"00",X"01",X"FE",X"1D",X"00",X"00",X"29",
		X"00",X"00",X"2A",X"01",X"FC",X"1D",X"39",X"3A",
		X"FC",X"FF",X"21",X"21",X"28",X"51",X"29",X"1A",
		X"02",X"16",X"2A",X"17",X"1B",X"03",X"CB",X"E2",
		X"01",X"49",X"01",X"00",X"67",X"26",X"03",X"CB",
		X"F0",X"24",X"01",X"00",X"26",X"03",X"CB",X"E3",
		X"28",X"66",X"01",X"28",X"24",X"25",X"00",X"29",
		X"2A",X"00",X"29",X"01",X"29",X"6A",X"03",X"04",
		X"68",X"01",X"CB",X"EF",X"4D",X"61",X"6E",X"64",
		X"65",X"6C",X"62",X"72",X"20",X"18",X"54",X"FB",
		X"EE",X"19",X"02",X"00",X"DF",X"11",X"01",X"01",
		X"2B",X"30",X"CD",X"CE",X"11",X"A7",X"04",X"2B",
		X"22",X"B4",X"FD",X"2B",X"32",X"1A",X"33",X"E6",
		X"78",X"35",X"53",X"05",X"E3",X"80",X"5E",X"33",
		X"21",X"32",X"2B",X"34",X"E3",X"40",X"5E",X"34",
		X"59",X"00",X"2B",X"36",X"2B",X"38",X"21",X"38",
		X"35",X"4D",X"5F",X"21",X"36",X"35",X"72",X"5D",
		X"21",X"3A",X"7F",X"00",X"5E",X"24",X"21",X"3A",
		X"7F",X"01",X"5E",X"25",X"21",X"3A",X"7F",X"02",
		X"5E",X"26",X"21",X"3A",X"E3",X"03",X"2B",X"3A",
		X"82",X"FF",X"8C",X"F9",X"35",X"72",X"56",X"21",
		X"3A",X"E3",X"07",X"2B",X"3A",X"11",X"C0",X"06",
		X"2B",X"22",X"B4",X"F2",X"21",X"38",X"35",X"53",
		X"77",X"59",X"24",X"99",X"36",X"AD",X"2B",X"38",
		X"35",X"72",X"6D",X"FF",X"21",X"36",X"E3",X"01",
		X"82",X"03",X"2B",X"36",X"90",X"A5",X"35",X"56",
		X"88",X"59",X"3F",X"00",X"FD",X"04",X"68",X"18",
		X"F0",X"32",X"21",X"38",X"E6",X"01",X"2B",X"38",
		X"93",X"32",X"90",X"A5",X"59",X"24",X"99",X"36",
		X"AD",X"35",X"3F",X"98",X"8C",X"3F",X"F0",X"32",
		X"93",X"32",X"90",X"9D",X"11",X"FF",X"FF",X"2B",
		X"38",X"21",X"36",X"E3",X"01",X"82",X"03",X"2B",
		X"36",X"21",X"32",X"B8",X"34",X"35",X"72",X"C8",
		X"59",X"00",X"F0",X"32",X"21",X"32",X"E6",X"40",
		X"5E",X"32",X"93",X"33",X"21",X"32",X"35",X"53",
		X"C4",X"11",X"00",X"88",X"99",X"32",X"2B",X"32",
		X"1A",X"33",X"5E",X"35",X"1A",X"0E",X"F0",X"30",
		X"90",X"27",X"2B",X"3C",X"11",X"00",X"13",X"2B",
		X"3A",X"CF",X"3C",X"CF",X"3C",X"CF",X"3C",X"90",
		X"D0",X"00",X"50",X"69",X"63",X"74",X"75",X"72",
		X"65",X"73",X"7A",X"18",X"59",X"FB",X"EE",X"19",
		X"02",X"00",X"95",X"CD",X"43",X"E6",X"52",X"35",
		X"53",X"0E",X"E3",X"32",X"2B",X"30",X"11",X"00",
		X"07",X"90",X"13",X"2B",X"30",X"11",X"00",X"08",
		X"2B",X"32",X"21",X"30",X"E9",X"E9",X"99",X"30",
		X"99",X"32",X"2B",X"32",X"21",X"34",X"2B",X"28",
		X"E3",X"06",X"2B",X"34",X"59",X"05",X"2B",X"30",
		X"21",X"32",X"7F",X"00",X"5E",X"26",X"B4",X"CB",
		X"93",X"32",X"93",X"28",X"21",X"30",X"E6",X"01",
		X"35",X"4D",X"29",X"5E",X"26",X"B4",X"CB",X"FF",
		X"2B",X"36",X"11",X"E1",X"04",X"2B",X"22",X"11",
		X"20",X"0F",X"2B",X"24",X"11",X"06",X"50",X"2B",
		X"34",X"CD",X"65",X"20",X"52",X"65",X"61",X"64",
		X"79",X"20",X"74",X"6F",X"20",X"6C",X"6F",X"61",
		X"64",X"00",X"2B",X"38",X"21",X"38",X"AD",X"35",
		X"3F",X"73",X"93",X"38",X"CF",X"36",X"90",X"67",
		X"5E",X"28",X"11",X"0C",X"59",X"2B",X"3A",X"11",
		X"0C",X"5B",X"2B",X"3C",X"59",X"67",X"5E",X"26",
		X"11",X"07",X"59",X"00",X"FD",X"04",X"68",X"18",
		X"2B",X"3E",X"11",X"58",X"59",X"2B",X"40",X"11",
		X"0C",X"5A",X"2B",X"1A",X"FF",X"5A",X"0C",X"75",
		X"21",X"3C",X"2B",X"24",X"59",X"CF",X"5E",X"27",
		X"21",X"3E",X"2B",X"22",X"B4",X"FE",X"59",X"DB",
		X"5E",X"27",X"B4",X"FE",X"59",X"EB",X"5E",X"27",
		X"B4",X"FE",X"59",X"FB",X"5E",X"27",X"B4",X"FE",
		X"21",X"40",X"2B",X"22",X"B4",X"FD",X"59",X"02",
		X"5E",X"27",X"21",X"3E",X"2B",X"22",X"B4",X"FE",
		X"59",X"06",X"5E",X"27",X"21",X"40",X"2B",X"22",
		X"B4",X"FD",X"21",X"3E",X"2B",X"22",X"B4",X"FE",
		X"1A",X"27",X"E3",X"04",X"5E",X"27",X"8C",X"F2",
		X"35",X"72",X"3E",X"59",X"B9",X"5E",X"27",X"B4",
		X"FE",X"1A",X"26",X"35",X"72",X"64",X"59",X"0C",
		X"90",X"66",X"59",X"03",X"F0",X"3A",X"1A",X"3A",
		X"E6",X"0B",X"82",X"7F",X"E3",X"0C",X"5E",X"3A",
		X"59",X"3F",X"F0",X"3A",X"11",X"1C",X"59",X"2B",
		X"22",X"B4",X"EE",X"90",X"0A",X"00",X"4C",X"6F",
		X"61",X"64",X"65",X"72",X"00",X"00",X"70",X"18",
		X"5A",X"FB",X"EE",X"19",X"02",X"00",X"D4",X"CD",
		X"25",X"75",X"21",X"30",X"AD",X"2B",X"32",X"35",
		X"3F",X"23",X"93",X"30",X"21",X"32",X"8C",X"0A",
		X"35",X"72",X"1F",X"59",X"02",X"5E",X"34",X"11",
		X"00",X"08",X"99",X"34",X"2B",X"34",X"90",X"21",
		X"CF",X"36",X"90",X"01",X"63",X"FF",X"2B",X"38",
		X"CD",X"CD",X"54",X"68",X"69",X"73",X"20",X"47",
		X"69",X"67",X"61",X"74",X"72",X"6F",X"6E",X"20",
		X"54",X"54",X"4C",X"20",X"63",X"6F",X"6D",X"70",
		X"75",X"74",X"65",X"72",X"0A",X"6B",X"69",X"74",
		X"20",X"77",X"61",X"73",X"20",X"62",X"72",X"6F",
		X"75",X"67",X"68",X"74",X"20",X"74",X"6F",X"20",
		X"79",X"6F",X"75",X"20",X"62",X"79",X"0A",X"4D",
		X"61",X"72",X"63",X"00",X"FD",X"04",X"68",X"18",
		X"65",X"6C",X"20",X"76",X"61",X"6E",X"20",X"4B",
		X"65",X"72",X"76",X"69",X"6E",X"63",X"6B",X"20",
		X"61",X"6E",X"64",X"0A",X"57",X"61",X"6C",X"74",
		X"65",X"72",X"20",X"42",X"65",X"6C",X"67",X"65",
		X"72",X"73",X"2E",X"0A",X"0A",X"60",X"54",X"65",
		X"74",X"72",X"6F",X"6E",X"69",X"73",X"27",X"20",
		X"69",X"73",X"20",X"62",X"79",X"20",X"61",X"74",
		X"36",X"37",X"20",X"61",X"6E",X"64",X"0A",X"60",
		X"42",X"72",X"69",X"63",X"6B",X"73",X"27",X"20",
		X"62",X"79",X"20",X"78",X"62",X"78",X"2E",X"0A",
		X"0A",X"53",X"70",X"65",X"63",X"69",X"61",X"6C",
		X"20",X"74",X"68",X"61",X"6E",X"6B",X"73",X"20",
		X"6D",X"75",X"73",X"74",X"20",X"67",X"6F",X"20",
		X"74",X"6F",X"00",X"2B",X"3A",X"93",X"1B",X"FF",
		X"03",X"00",X"E8",X"CD",X"98",X"0A",X"4D",X"61",
		X"72",X"63",X"2C",X"20",X"50",X"61",X"75",X"6C",
		X"2C",X"20",X"49",X"76",X"61",X"6E",X"61",X"2C",
		X"20",X"4F",X"73",X"63",X"61",X"72",X"2C",X"0A",
		X"4D",X"61",X"72",X"74",X"69",X"6A",X"6E",X"2C",
		X"20",X"45",X"72",X"69",X"6B",X"2C",X"20",X"43",
		X"68",X"75",X"63",X"6B",X"2C",X"20",X"42",X"65",
		X"6E",X"2C",X"0A",X"44",X"69",X"65",X"74",X"65",
		X"72",X"2C",X"20",X"4D",X"61",X"72",X"74",X"69",
		X"6E",X"2C",X"20",X"42",X"72",X"61",X"64",X"2C",
		X"20",X"4C",X"6F",X"75",X"2C",X"0A",X"50",X"68",
		X"69",X"6C",X"2C",X"20",X"42",X"72",X"69",X"61",
		X"6E",X"2C",X"20",X"44",X"61",X"76",X"69",X"64",
		X"2C",X"20",X"44",X"61",X"76",X"65",X"2C",X"0A",
		X"48",X"47",X"20",X"61",X"6E",X"64",X"20",X"61",
		X"6C",X"6C",X"20",X"66",X"61",X"6E",X"73",X"21",
		X"0A",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"00",X"FD",X"04",X"68",X"18",
		X"20",X"4D",X"61",X"72",X"63",X"65",X"6C",X"20",
		X"26",X"20",X"57",X"61",X"6C",X"74",X"65",X"72",
		X"0A",X"00",X"2B",X"3C",X"CD",X"CD",X"11",X"00",
		X"08",X"2B",X"3E",X"11",X"01",X"88",X"2B",X"40",
		X"59",X"00",X"5E",X"24",X"5E",X"25",X"11",X"E1",
		X"04",X"2B",X"22",X"21",X"3E",X"2B",X"28",X"B4",
		X"CB",X"11",X"00",X"08",X"99",X"3E",X"2B",X"3E",
		X"35",X"4D",X"B3",X"99",X"40",X"2B",X"3E",X"82",
		X"FF",X"8C",X"A0",X"35",X"72",X"B1",X"FF",X"2B",
		X"42",X"CD",X"E1",X"1A",X"0E",X"99",X"44",X"82",
		X"FF",X"2B",X"46",X"1A",X"0E",X"B8",X"46",X"35",
		X"72",X"D9",X"FF",X"2B",X"48",X"93",X"1B",X"FF",
		X"04",X"00",X"81",X"CD",X"4A",X"21",X"32",X"E6",
		X"52",X"35",X"53",X"10",X"E3",X"32",X"2B",X"40",
		X"11",X"00",X"07",X"90",X"15",X"2B",X"40",X"11",
		X"00",X"08",X"2B",X"4A",X"21",X"40",X"E9",X"E9",
		X"99",X"40",X"99",X"4A",X"2B",X"4A",X"21",X"4C",
		X"5E",X"25",X"21",X"34",X"2B",X"28",X"E3",X"06",
		X"2B",X"34",X"11",X"E1",X"04",X"2B",X"22",X"59",
		X"FB",X"2B",X"40",X"21",X"4A",X"7F",X"00",X"93",
		X"4A",X"5E",X"26",X"B4",X"CB",X"93",X"28",X"93",
		X"40",X"21",X"40",X"35",X"72",X"36",X"FF",X"2B",
		X"36",X"11",X"02",X"08",X"2B",X"34",X"CF",X"42",
		X"59",X"3E",X"2B",X"4C",X"11",X"00",X"08",X"2B",
		X"34",X"21",X"3A",X"2B",X"30",X"CF",X"38",X"21",
		X"3C",X"2B",X"30",X"CF",X"38",X"59",X"F0",X"2B",
		X"44",X"CF",X"48",X"21",X"4C",X"8C",X"08",X"35",
		X"3F",X"7D",X"21",X"4C",X"E6",X"09",X"2B",X"4C",
		X"90",X"57",X"90",X"53",X"00",X"43",X"72",X"65",
		X"64",X"69",X"74",X"73",X"00",X"94",X"18",X"5B",
		X"FB",X"EE",X"19",X"00",X"4A",X"4E",X"A1",X"2D",
		X"A1",X"21",X"A1",X"00",X"FD",X"04",X"68",X"18",
		X"19",X"A1",X"1E",X"00",X"03",X"00",X"06",X"B6",
		X"2D",X"A1",X"22",X"A1",X"15",X"A1",X"2B",X"A1",
		X"2A",X"A1",X"1B",X"A1",X"16",X"A1",X"2E",X"D5",
		X"30",X"A1",X"30",X"00",X"05",X"A1",X"28",X"A1",
		X"2C",X"A1",X"26",X"A1",X"25",X"A1",X"29",X"00",
		X"04",X"A1",X"1A",X"C7",X"23",X"A1",X"1F",X"A1",
		X"24",X"01",X"00",X"A1",X"23",X"A1",X"20",X"E4",
		X"1C",X"A1",X"1D",X"CC",X"1C",X"A1",X"1C",X"CC",
		X"1D",X"A1",X"18",X"C2",X"16",X"A1",X"17",X"A1",
		X"2F",X"02",X"00",X"F4",X"11",X"00",X"08",X"2B",
		X"CE",X"11",X"00",X"07",X"2B",X"D2",X"11",X"A1",
		X"7A",X"2B",X"D4",X"11",X"01",X"01",X"2B",X"D0",
		X"CF",X"64",X"CF",X"62",X"CF",X"60",X"CF",X"5E",
		X"CF",X"5C",X"CF",X"5A",X"11",X"00",X"00",X"2B",
		X"DE",X"2B",X"E0",X"2B",X"C2",X"11",X"32",X"00",
		X"2B",X"C8",X"2B",X"C6",X"1A",X"06",X"5E",X"38",
		X"59",X"00",X"5E",X"37",X"1A",X"0E",X"2B",X"C4",
		X"11",X"E0",X"08",X"2B",X"BA",X"CF",X"58",X"1A",
		X"0E",X"5E",X"40",X"5E",X"CC",X"CF",X"56",X"CF",
		X"54",X"CF",X"96",X"CF",X"52",X"5E",X"36",X"8C",
		X"FB",X"35",X"3F",X"5F",X"1A",X"36",X"35",X"72",
		X"6E",X"21",X"C8",X"2B",X"C6",X"21",X"C2",X"E3",
		X"01",X"2B",X"C2",X"B8",X"C6",X"35",X"50",X"49",
		X"59",X"00",X"5E",X"36",X"1A",X"37",X"35",X"72",
		X"75",X"CF",X"50",X"21",X"A4",X"99",X"AC",X"35",
		X"53",X"85",X"11",X"00",X"00",X"B8",X"AC",X"2B",
		X"A4",X"90",X"99",X"21",X"A4",X"99",X"A8",X"99",
		X"AC",X"E6",X"0A",X"35",X"56",X"99",X"11",X"0A",
		X"00",X"B8",X"A8",X"B8",X"AC",X"2B",X"A4",X"21",
		X"C2",X"B8",X"C6",X"35",X"50",X"C4",X"11",X"00",
		X"00",X"2B",X"C2",X"59",X"00",X"5E",X"37",X"93",
		X"A6",X"21",X"A6",X"00",X"FD",X"04",X"68",X"18",
		X"99",X"AA",X"E6",X"14",X"35",X"56",X"C4",X"1A",
		X"A6",X"E6",X"01",X"5E",X"A6",X"CF",X"4E",X"CF",
		X"58",X"59",X"FF",X"5E",X"37",X"90",X"45",X"CF",
		X"4C",X"21",X"C0",X"35",X"3F",X"EE",X"E6",X"01",
		X"35",X"72",X"D9",X"CF",X"64",X"11",X"A1",X"34",
		X"2B",X"3A",X"90",X"18",X"1A",X"36",X"35",X"3F",
		X"E2",X"CF",X"4A",X"90",X"EE",X"1A",X"A6",X"E6",
		X"01",X"5E",X"A6",X"CF",X"4E",X"CF",X"58",X"90",
		X"45",X"CF",X"4E",X"90",X"45",X"03",X"00",X"71",
		X"1A",X"11",X"8C",X"FF",X"35",X"72",X"08",X"5E",
		X"35",X"FF",X"1A",X"11",X"8C",X"FB",X"35",X"72",
		X"17",X"11",X"02",X"00",X"2B",X"C6",X"1A",X"11",
		X"FF",X"1A",X"35",X"35",X"3F",X"1F",X"1A",X"00",
		X"FF",X"1A",X"11",X"5E",X"35",X"8C",X"FD",X"35",
		X"72",X"31",X"21",X"A4",X"E6",X"01",X"2B",X"A4",
		X"1A",X"11",X"FF",X"1A",X"11",X"8C",X"FE",X"35",
		X"72",X"41",X"21",X"A4",X"E3",X"01",X"2B",X"A4",
		X"1A",X"11",X"FF",X"1A",X"11",X"8C",X"F7",X"35",
		X"72",X"6C",X"21",X"9E",X"2B",X"CC",X"E3",X"10",
		X"82",X"30",X"2B",X"9E",X"75",X"CF",X"82",X"63",
		X"21",X"A6",X"99",X"AA",X"99",X"AE",X"E6",X"14",
		X"35",X"56",X"6C",X"21",X"CC",X"2B",X"9E",X"75",
		X"CF",X"82",X"63",X"1A",X"00",X"FF",X"1A",X"11",
		X"FF",X"04",X"00",X"96",X"11",X"A1",X"0F",X"2B",
		X"CC",X"21",X"DC",X"E6",X"01",X"99",X"CC",X"AD",
		X"2B",X"E4",X"1A",X"E0",X"E3",X"01",X"5E",X"9A",
		X"11",X"00",X"00",X"2B",X"CC",X"21",X"CC",X"99",
		X"E4",X"2B",X"CC",X"1A",X"9A",X"E6",X"01",X"5E",
		X"9A",X"35",X"72",X"17",X"21",X"CC",X"2B",X"E4",
		X"99",X"DE",X"2B",X"DE",X"11",X"A6",X"0F",X"2B",
		X"CC",X"21",X"E0",X"E9",X"99",X"CC",X"F6",X"B8",
		X"DE",X"35",X"4D",X"00",X"FD",X"04",X"68",X"18",
		X"78",X"2B",X"DE",X"11",X"00",X"00",X"B8",X"DE",
		X"2B",X"DE",X"1A",X"E0",X"8C",X"08",X"35",X"3F",
		X"78",X"21",X"C8",X"E6",X"05",X"2B",X"C8",X"2B",
		X"C6",X"93",X"E0",X"75",X"CF",X"6E",X"63",X"11",
		X"AF",X"7F",X"2B",X"D6",X"11",X"5F",X"6D",X"2B",
		X"D8",X"75",X"CF",X"6C",X"63",X"11",X"B2",X"7F",
		X"2B",X"D6",X"11",X"3A",X"6D",X"2B",X"D8",X"75",
		X"CF",X"6C",X"63",X"75",X"CF",X"6A",X"63",X"11",
		X"A1",X"7F",X"2B",X"D6",X"11",X"44",X"6D",X"2B",
		X"D8",X"75",X"CF",X"6C",X"63",X"21",X"E4",X"E6",
		X"05",X"2B",X"E4",X"35",X"4D",X"78",X"FF",X"05",
		X"00",X"8C",X"11",X"A7",X"7F",X"2B",X"CC",X"AD",
		X"E3",X"05",X"5E",X"9A",X"8C",X"3A",X"35",X"3F",
		X"12",X"1A",X"9A",X"F0",X"CC",X"FF",X"59",X"30",
		X"F0",X"CC",X"11",X"A6",X"7F",X"2B",X"CC",X"AD",
		X"E3",X"01",X"5E",X"9A",X"8C",X"3A",X"35",X"3F",
		X"2A",X"1A",X"9A",X"F0",X"CC",X"FF",X"59",X"30",
		X"F0",X"CC",X"11",X"A5",X"7F",X"2B",X"CC",X"AD",
		X"E3",X"01",X"5E",X"9A",X"8C",X"3A",X"35",X"3F",
		X"42",X"1A",X"9A",X"F0",X"CC",X"FF",X"59",X"30",
		X"F0",X"CC",X"11",X"A4",X"7F",X"2B",X"CC",X"AD",
		X"E3",X"01",X"5E",X"9A",X"8C",X"3A",X"35",X"3F",
		X"5A",X"1A",X"9A",X"F0",X"CC",X"FF",X"59",X"30",
		X"F0",X"CC",X"11",X"A3",X"7F",X"2B",X"CC",X"AD",
		X"E3",X"01",X"5E",X"9A",X"8C",X"3A",X"35",X"3F",
		X"72",X"1A",X"9A",X"F0",X"CC",X"FF",X"59",X"30",
		X"F0",X"CC",X"11",X"A2",X"7F",X"2B",X"CC",X"AD",
		X"E3",X"01",X"5E",X"9A",X"8C",X"3A",X"35",X"3F",
		X"89",X"1A",X"9A",X"F0",X"CC",X"FF",X"06",X"00",
		X"0C",X"1A",X"0E",X"B8",X"C4",X"35",X"3F",X"FE",
		X"1A",X"0E",X"2B",X"C4",X"FF",X"08",X"A1",X"40",
		X"3C",X"3C",X"04",X"00",X"FD",X"04",X"68",X"18",
		X"01",X"00",X"01",X"00",X"01",X"01",X"01",X"02",
		X"01",X"03",X"01",X"00",X"00",X"3C",X"3C",X"01",
		X"04",X"02",X"00",X"02",X"00",X"02",X"01",X"02",
		X"02",X"02",X"03",X"00",X"00",X"3C",X"3C",X"04",
		X"01",X"00",X"02",X"00",X"02",X"01",X"02",X"02",
		X"02",X"03",X"02",X"00",X"00",X"3C",X"3C",X"01",
		X"04",X"01",X"00",X"01",X"00",X"01",X"01",X"01",
		X"02",X"01",X"03",X"00",X"00",X"08",X"E0",X"10",
		X"A1",X"08",X"A1",X"09",X"A1",X"0A",X"A1",X"0B",
		X"A1",X"0C",X"A1",X"0D",X"A1",X"0E",X"A1",X"08",
		X"09",X"A1",X"40",X"30",X"30",X"03",X"02",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"02",
		X"01",X"00",X"00",X"30",X"30",X"02",X"03",X"01",
		X"00",X"01",X"00",X"02",X"00",X"01",X"01",X"01",
		X"02",X"00",X"00",X"30",X"30",X"03",X"02",X"00",
		X"01",X"00",X"01",X"01",X"01",X"02",X"01",X"02",
		X"02",X"00",X"00",X"30",X"30",X"02",X"03",X"00",
		X"00",X"01",X"00",X"01",X"01",X"00",X"02",X"01",
		X"02",X"00",X"00",X"0A",X"A1",X"40",X"0B",X"0B",
		X"03",X"02",X"00",X"00",X"02",X"00",X"00",X"01",
		X"01",X"01",X"02",X"01",X"00",X"00",X"0B",X"0B",
		X"02",X"03",X"01",X"00",X"01",X"00",X"01",X"01",
		X"01",X"02",X"02",X"02",X"00",X"00",X"0B",X"0B",
		X"03",X"02",X"00",X"01",X"00",X"01",X"01",X"01",
		X"02",X"01",X"00",X"02",X"00",X"00",X"0B",X"0B",
		X"02",X"03",X"00",X"00",X"00",X"00",X"01",X"00",
		X"01",X"01",X"01",X"02",X"00",X"00",X"0B",X"A1",
		X"40",X"0F",X"0F",X"02",X"02",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"01",X"01",X"01",X"00",
		X"00",X"0F",X"0F",X"02",X"02",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"01",X"01",X"01",X"00",
		X"00",X"0F",X"0F",X"00",X"FD",X"04",X"68",X"18",
		X"02",X"02",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"01",X"01",X"01",X"00",X"00",X"0F",X"0F",
		X"02",X"02",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"01",X"01",X"01",X"00",X"00",X"0C",X"A1",
		X"40",X"0C",X"0C",X"03",X"02",X"00",X"00",X"01",
		X"00",X"02",X"00",X"00",X"01",X"01",X"01",X"00",
		X"00",X"0C",X"0C",X"02",X"03",X"01",X"00",X"01",
		X"00",X"01",X"01",X"02",X"01",X"02",X"02",X"00",
		X"00",X"0C",X"0C",X"03",X"02",X"00",X"01",X"01",
		X"01",X"02",X"01",X"00",X"02",X"01",X"02",X"00",
		X"00",X"0C",X"0C",X"02",X"03",X"00",X"00",X"00",
		X"00",X"00",X"01",X"01",X"01",X"01",X"02",X"00",
		X"00",X"0D",X"A1",X"40",X"33",X"33",X"03",X"02",
		X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"01",
		X"02",X"01",X"00",X"00",X"33",X"33",X"02",X"03",
		X"01",X"00",X"01",X"00",X"01",X"01",X"02",X"01",
		X"01",X"02",X"00",X"00",X"33",X"33",X"03",X"02",
		X"00",X"01",X"00",X"01",X"01",X"01",X"02",X"01",
		X"01",X"02",X"00",X"00",X"33",X"33",X"02",X"03",
		X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"01",
		X"01",X"02",X"00",X"00",X"0E",X"A1",X"40",X"03",
		X"03",X"03",X"02",X"00",X"00",X"00",X"00",X"01",
		X"00",X"01",X"01",X"02",X"01",X"00",X"00",X"03",
		X"03",X"02",X"03",X"01",X"00",X"02",X"00",X"01",
		X"01",X"02",X"01",X"01",X"02",X"00",X"00",X"03",
		X"03",X"03",X"02",X"00",X"01",X"00",X"01",X"01",
		X"01",X"01",X"02",X"02",X"02",X"00",X"00",X"03",
		X"03",X"02",X"03",X"00",X"00",X"01",X"00",X"00",
		X"01",X"01",X"01",X"00",X"02",X"00",X"00",X"0F",
		X"A1",X"04",X"0A",X"19",X"32",X"64",X"0F",X"A6",
		X"12",X"FA",X"00",X"EE",X"02",X"E8",X"03",X"D0",
		X"07",X"A0",X"0F",X"00",X"FD",X"04",X"68",X"18",
		X"40",X"1F",X"80",X"3E",X"00",X"7D",X"00",X"FA",
		X"15",X"A1",X"4F",X"11",X"D4",X"04",X"2B",X"22",
		X"11",X"00",X"00",X"2B",X"24",X"2B",X"26",X"59",
		X"14",X"5E",X"99",X"59",X"3C",X"5E",X"98",X"59",
		X"50",X"5E",X"9B",X"59",X"0A",X"5E",X"9A",X"21",
		X"CE",X"99",X"98",X"2B",X"28",X"B4",X"FF",X"1A",
		X"98",X"E3",X"04",X"5E",X"98",X"1A",X"9A",X"E6",
		X"01",X"5E",X"9A",X"35",X"72",X"BB",X"1A",X"99",
		X"E3",X"01",X"5E",X"99",X"59",X"3C",X"5E",X"98",
		X"75",X"CF",X"96",X"63",X"59",X"0A",X"5E",X"9A",
		X"1A",X"9B",X"E6",X"01",X"5E",X"9B",X"35",X"72",
		X"BB",X"FF",X"16",X"A1",X"32",X"11",X"D4",X"04",
		X"2B",X"22",X"11",X"00",X"00",X"2B",X"24",X"2B",
		X"26",X"59",X"3C",X"5E",X"9B",X"59",X"28",X"5E",
		X"9A",X"11",X"00",X"08",X"2B",X"98",X"11",X"00",
		X"7F",X"2B",X"30",X"75",X"CF",X"94",X"2B",X"CC",
		X"59",X"00",X"F0",X"CC",X"21",X"CC",X"E3",X"5F",
		X"2B",X"CC",X"59",X"00",X"F0",X"CC",X"FF",X"17",
		X"A1",X"4A",X"63",X"21",X"98",X"2B",X"28",X"B4",
		X"FF",X"21",X"30",X"2B",X"28",X"B4",X"FF",X"1A",
		X"98",X"E3",X"04",X"5E",X"98",X"1A",X"30",X"E3",
		X"04",X"5E",X"30",X"1A",X"9A",X"E6",X"01",X"5E",
		X"9A",X"35",X"72",X"A0",X"75",X"21",X"98",X"CF",
		X"92",X"63",X"75",X"21",X"30",X"CF",X"92",X"63",
		X"93",X"99",X"1A",X"31",X"E6",X"01",X"5E",X"31",
		X"59",X"00",X"5E",X"98",X"5E",X"30",X"59",X"28",
		X"5E",X"9A",X"1A",X"9B",X"E6",X"01",X"5E",X"9B",
		X"35",X"72",X"A0",X"FF",X"18",X"A1",X"3B",X"11",
		X"D4",X"04",X"2B",X"22",X"21",X"BE",X"2B",X"24",
		X"2B",X"26",X"59",X"04",X"5E",X"9B",X"1A",X"98",
		X"E9",X"E9",X"E3",X"3C",X"5E",X"98",X"1A",X"99",
		X"E9",X"E9",X"E3",X"00",X"FD",X"04",X"68",X"18",
		X"14",X"5E",X"99",X"21",X"CE",X"99",X"98",X"2B",
		X"28",X"B4",X"FF",X"75",X"CF",X"96",X"63",X"1A",
		X"99",X"E3",X"01",X"5E",X"99",X"1A",X"9B",X"E6",
		X"01",X"5E",X"9B",X"35",X"72",X"BE",X"FF",X"19",
		X"A1",X"4C",X"21",X"9C",X"99",X"BA",X"F6",X"99",
		X"9E",X"2B",X"BC",X"F6",X"2B",X"BE",X"21",X"BC",
		X"E3",X"05",X"2B",X"BC",X"59",X"04",X"5E",X"9A",
		X"21",X"BC",X"E3",X"01",X"2B",X"BC",X"AD",X"99",
		X"A4",X"5E",X"98",X"35",X"50",X"E1",X"E6",X"0A",
		X"35",X"53",X"E1",X"21",X"BC",X"E3",X"01",X"2B",
		X"BC",X"AD",X"99",X"A6",X"B8",X"AE",X"5E",X"99",
		X"35",X"50",X"E1",X"E6",X"14",X"35",X"53",X"E1",
		X"75",X"CF",X"90",X"63",X"1A",X"9A",X"E6",X"01",
		X"5E",X"9A",X"35",X"72",X"B5",X"FF",X"1A",X"A1",
		X"5D",X"21",X"A0",X"99",X"BA",X"F6",X"99",X"A2",
		X"2B",X"BC",X"F6",X"2B",X"BE",X"21",X"BC",X"E3",
		X"02",X"F6",X"2B",X"30",X"21",X"BC",X"E3",X"04",
		X"F6",X"2B",X"32",X"21",X"BC",X"E3",X"05",X"2B",
		X"BC",X"59",X"04",X"5E",X"9A",X"11",X"61",X"17",
		X"2B",X"98",X"75",X"CF",X"8E",X"63",X"1A",X"98",
		X"2B",X"CC",X"21",X"BC",X"E3",X"01",X"2B",X"BC",
		X"AD",X"99",X"CC",X"5E",X"98",X"1A",X"99",X"2B",
		X"CC",X"21",X"BC",X"E3",X"01",X"2B",X"BC",X"AD",
		X"99",X"CC",X"5E",X"99",X"21",X"BE",X"F0",X"98",
		X"75",X"CF",X"96",X"63",X"1A",X"9A",X"E6",X"01",
		X"5E",X"9A",X"35",X"72",X"C3",X"FF",X"1B",X"A1",
		X"56",X"11",X"15",X"15",X"2B",X"BE",X"75",X"CF",
		X"8C",X"63",X"11",X"FF",X"00",X"2B",X"A6",X"11",
		X"FF",X"00",X"2B",X"A4",X"59",X"0C",X"5E",X"9A",
		X"75",X"CF",X"8A",X"63",X"11",X"14",X"00",X"2B",
		X"A6",X"11",X"FF",X"00",X"2B",X"A4",X"59",X"0C",
		X"5E",X"9A",X"75",X"00",X"FD",X"04",X"68",X"18",
		X"CF",X"8A",X"63",X"75",X"CF",X"88",X"63",X"11",
		X"FF",X"00",X"2B",X"A6",X"11",X"FF",X"00",X"2B",
		X"A4",X"59",X"15",X"5E",X"9A",X"75",X"CF",X"86",
		X"63",X"11",X"FF",X"00",X"2B",X"A6",X"11",X"0A",
		X"00",X"2B",X"A4",X"59",X"15",X"5E",X"9A",X"75",
		X"CF",X"86",X"63",X"FF",X"1C",X"A1",X"5B",X"11",
		X"38",X"15",X"2B",X"98",X"11",X"38",X"16",X"2B",
		X"30",X"11",X"38",X"17",X"2B",X"32",X"59",X"30",
		X"5E",X"9A",X"59",X"15",X"F0",X"98",X"F0",X"30",
		X"F0",X"32",X"93",X"98",X"93",X"30",X"93",X"32",
		X"1A",X"9A",X"E6",X"01",X"5E",X"9A",X"35",X"72",
		X"B2",X"FF",X"21",X"A6",X"5E",X"99",X"21",X"A4",
		X"5E",X"98",X"75",X"CF",X"90",X"63",X"93",X"A4",
		X"1A",X"9A",X"E6",X"01",X"5E",X"9A",X"35",X"72",
		X"CA",X"FF",X"21",X"A6",X"5E",X"99",X"21",X"A4",
		X"5E",X"98",X"75",X"CF",X"90",X"63",X"93",X"A6",
		X"1A",X"9A",X"E6",X"01",X"5E",X"9A",X"35",X"72",
		X"E2",X"FF",X"1D",X"A1",X"44",X"11",X"38",X"70",
		X"2B",X"98",X"11",X"38",X"71",X"2B",X"30",X"11",
		X"38",X"72",X"2B",X"32",X"59",X"30",X"5E",X"9A",
		X"59",X"15",X"F0",X"98",X"F0",X"30",X"F0",X"32",
		X"93",X"98",X"93",X"30",X"93",X"32",X"1A",X"9A",
		X"E6",X"01",X"5E",X"9A",X"35",X"72",X"B2",X"FF",
		X"21",X"30",X"B8",X"32",X"2B",X"CC",X"1A",X"CC",
		X"8C",X"02",X"35",X"72",X"D9",X"93",X"98",X"1A",
		X"CD",X"8C",X"02",X"35",X"72",X"E2",X"93",X"99",
		X"FF",X"1E",X"A1",X"4E",X"21",X"B6",X"99",X"BA",
		X"F6",X"99",X"B8",X"2B",X"BC",X"11",X"00",X"00",
		X"2B",X"BE",X"21",X"BC",X"E3",X"05",X"2B",X"BC",
		X"59",X"04",X"5E",X"9A",X"21",X"BC",X"E3",X"01",
		X"2B",X"BC",X"AD",X"99",X"B0",X"5E",X"98",X"35",
		X"50",X"E3",X"E6",X"00",X"FD",X"04",X"68",X"18",
		X"0A",X"35",X"53",X"E3",X"21",X"BC",X"E3",X"01",
		X"2B",X"BC",X"AD",X"99",X"B2",X"B8",X"B4",X"5E",
		X"99",X"35",X"50",X"E3",X"E6",X"14",X"35",X"53",
		X"E3",X"75",X"CF",X"90",X"63",X"1A",X"9A",X"E6",
		X"01",X"5E",X"9A",X"35",X"72",X"B7",X"FF",X"1F",
		X"A1",X"3E",X"11",X"D4",X"04",X"2B",X"22",X"11",
		X"15",X"15",X"2B",X"24",X"2B",X"26",X"59",X"06",
		X"5E",X"9A",X"59",X"62",X"5E",X"28",X"59",X"16",
		X"5E",X"29",X"B4",X"FF",X"21",X"28",X"E6",X"01",
		X"2B",X"CC",X"59",X"15",X"F0",X"CC",X"21",X"CC",
		X"E6",X"01",X"2B",X"CC",X"59",X"15",X"F0",X"CC",
		X"1A",X"29",X"E3",X"01",X"5E",X"29",X"1A",X"9A",
		X"E6",X"01",X"5E",X"9A",X"35",X"72",X"B7",X"FF",
		X"20",X"A1",X"1C",X"1A",X"98",X"E9",X"E9",X"E3",
		X"3C",X"5E",X"98",X"1A",X"99",X"E9",X"E9",X"E3",
		X"14",X"5E",X"99",X"21",X"CE",X"99",X"98",X"AD",
		X"2B",X"C0",X"75",X"CF",X"96",X"63",X"FF",X"21",
		X"A1",X"5E",X"21",X"9C",X"99",X"BA",X"F6",X"99",
		X"9E",X"2B",X"BC",X"E3",X"05",X"2B",X"BC",X"11",
		X"00",X"00",X"2B",X"C0",X"59",X"04",X"5E",X"9A",
		X"21",X"BC",X"E3",X"01",X"2B",X"BC",X"AD",X"99",
		X"A4",X"5E",X"98",X"35",X"50",X"F3",X"E6",X"0A",
		X"35",X"53",X"F3",X"21",X"BC",X"E3",X"01",X"2B",
		X"BC",X"AD",X"99",X"A6",X"B8",X"AE",X"5E",X"99",
		X"35",X"50",X"F3",X"E6",X"14",X"35",X"53",X"F3",
		X"75",X"CF",X"84",X"63",X"21",X"C0",X"35",X"3F",
		X"F3",X"21",X"A6",X"B8",X"AE",X"35",X"72",X"F2",
		X"11",X"01",X"00",X"2B",X"C0",X"FF",X"1A",X"9A",
		X"E6",X"01",X"5E",X"9A",X"35",X"72",X"B5",X"FF",
		X"22",X"A1",X"59",X"1A",X"38",X"82",X"07",X"E9",
		X"2B",X"9C",X"1A",X"38",X"82",X"30",X"2B",X"9E",
		X"75",X"CF",X"82",X"00",X"FD",X"04",X"68",X"18",
		X"63",X"11",X"FF",X"00",X"2B",X"A6",X"11",X"0A",
		X"00",X"B8",X"A8",X"E6",X"01",X"2B",X"CC",X"1A",
		X"07",X"82",X"07",X"E3",X"01",X"2B",X"CA",X"B8",
		X"CC",X"2B",X"CC",X"35",X"56",X"D3",X"21",X"CA",
		X"B8",X"CC",X"2B",X"CA",X"21",X"CA",X"B8",X"AC",
		X"2B",X"A4",X"75",X"CF",X"7E",X"63",X"75",X"CF",
		X"7C",X"63",X"75",X"CF",X"7A",X"63",X"75",X"CF",
		X"78",X"63",X"1A",X"DC",X"35",X"72",X"EF",X"FF",
		X"75",X"CF",X"76",X"63",X"75",X"CF",X"74",X"63",
		X"FF",X"23",X"A1",X"36",X"21",X"9C",X"99",X"BA",
		X"F6",X"99",X"9E",X"2B",X"BC",X"21",X"BC",X"E3",
		X"02",X"AD",X"2B",X"A8",X"21",X"BC",X"E3",X"03",
		X"AD",X"2B",X"AA",X"21",X"BC",X"E3",X"04",X"AD",
		X"2B",X"AC",X"21",X"BC",X"E3",X"05",X"AD",X"2B",
		X"AE",X"FF",X"1A",X"07",X"5E",X"38",X"82",X"07",
		X"E9",X"2B",X"A0",X"1A",X"38",X"82",X"30",X"2B",
		X"A2",X"FF",X"24",X"A1",X"44",X"59",X"03",X"5E",
		X"9A",X"11",X"00",X"00",X"2B",X"DC",X"59",X"13",
		X"5E",X"31",X"59",X"09",X"5E",X"30",X"21",X"30",
		X"2B",X"98",X"75",X"CF",X"84",X"63",X"21",X"C0",
		X"35",X"3F",X"CC",X"1A",X"30",X"E6",X"01",X"5E",
		X"30",X"35",X"53",X"B0",X"93",X"DC",X"75",X"CF",
		X"72",X"63",X"1A",X"31",X"E6",X"01",X"5E",X"31",
		X"35",X"53",X"AC",X"1A",X"9A",X"E6",X"01",X"5E",
		X"9A",X"35",X"53",X"A8",X"59",X"00",X"F0",X"D0",
		X"FF",X"25",X"A1",X"59",X"1A",X"31",X"5E",X"33",
		X"59",X"09",X"5E",X"32",X"1A",X"33",X"E6",X"01",
		X"5E",X"99",X"1A",X"32",X"5E",X"98",X"75",X"CF",
		X"84",X"63",X"1A",X"C0",X"5E",X"BE",X"5E",X"BF",
		X"21",X"32",X"2B",X"98",X"75",X"CF",X"90",X"63",
		X"1A",X"32",X"E6",X"01",X"5E",X"32",X"35",X"53",
		X"A7",X"75",X"CF",X"00",X"FD",X"04",X"68",X"18",
		X"70",X"63",X"1A",X"33",X"E6",X"01",X"5E",X"33",
		X"35",X"72",X"A3",X"59",X"09",X"5E",X"30",X"59",
		X"00",X"5E",X"99",X"1A",X"30",X"5E",X"98",X"11",
		X"00",X"00",X"2B",X"BE",X"75",X"CF",X"90",X"63",
		X"1A",X"30",X"E6",X"01",X"5E",X"30",X"35",X"53",
		X"DD",X"FF",X"26",X"A1",X"1B",X"1A",X"06",X"82",
		X"03",X"35",X"3F",X"B5",X"8C",X"01",X"35",X"3F",
		X"B0",X"59",X"00",X"F0",X"D0",X"FF",X"59",X"01",
		X"F0",X"D0",X"FF",X"59",X"FF",X"F0",X"D0",X"FF",
		X"27",X"A1",X"5D",X"11",X"E1",X"04",X"2B",X"22",
		X"59",X"00",X"5E",X"24",X"59",X"3F",X"5E",X"25",
		X"21",X"D6",X"AD",X"5E",X"34",X"93",X"D6",X"21",
		X"D6",X"AD",X"E6",X"20",X"2B",X"DA",X"2B",X"CC",
		X"E9",X"E9",X"99",X"DA",X"99",X"D2",X"2B",X"CC",
		X"21",X"DA",X"E6",X"32",X"35",X"50",X"D1",X"21",
		X"CC",X"E3",X"06",X"2B",X"CC",X"59",X"05",X"5E",
		X"9A",X"21",X"D8",X"2B",X"28",X"21",X"CC",X"7F",
		X"00",X"5E",X"26",X"B4",X"CB",X"93",X"CC",X"93",
		X"D8",X"1A",X"9A",X"E6",X"01",X"5E",X"9A",X"35",
		X"72",X"D5",X"93",X"D6",X"93",X"D8",X"1A",X"34",
		X"E6",X"01",X"5E",X"34",X"35",X"72",X"B3",X"FF",
		X"28",X"A1",X"5C",X"11",X"D4",X"04",X"2B",X"22",
		X"21",X"D6",X"AD",X"5E",X"34",X"93",X"D6",X"21",
		X"D6",X"AD",X"E6",X"30",X"2B",X"CC",X"E9",X"E9",
		X"99",X"D4",X"2B",X"CC",X"59",X"05",X"5E",X"9A",
		X"21",X"CC",X"F6",X"2B",X"24",X"21",X"CC",X"E3",
		X"02",X"AD",X"5E",X"26",X"59",X"15",X"5E",X"27",
		X"21",X"D8",X"2B",X"28",X"B4",X"FF",X"75",X"CF",
		X"96",X"63",X"93",X"CD",X"93",X"D9",X"1A",X"9A",
		X"E6",X"01",X"5E",X"9A",X"35",X"72",X"BC",X"93",
		X"D6",X"1A",X"D8",X"E3",X"04",X"5E",X"D8",X"1A",
		X"D9",X"E6",X"05",X"00",X"FD",X"04",X"68",X"18",
		X"5E",X"D9",X"1A",X"34",X"E6",X"01",X"5E",X"34",
		X"35",X"72",X"AB",X"FF",X"29",X"A1",X"5A",X"11",
		X"A9",X"7F",X"2B",X"E4",X"11",X"A2",X"7F",X"2B",
		X"CC",X"59",X"06",X"5E",X"9A",X"21",X"CC",X"AD",
		X"2B",X"E2",X"21",X"E4",X"AD",X"B8",X"E2",X"35",
		X"4D",X"F8",X"35",X"50",X"CA",X"93",X"E4",X"93",
		X"CC",X"1A",X"9A",X"E6",X"01",X"5E",X"9A",X"35",
		X"72",X"AD",X"11",X"A9",X"7F",X"2B",X"E4",X"11",
		X"A2",X"7F",X"2B",X"CC",X"59",X"06",X"5E",X"9A",
		X"21",X"CC",X"AD",X"F0",X"E4",X"93",X"E4",X"93",
		X"CC",X"1A",X"9A",X"E6",X"01",X"5E",X"9A",X"35",
		X"72",X"D8",X"11",X"A8",X"7F",X"2B",X"D6",X"11",
		X"44",X"16",X"2B",X"D8",X"75",X"CF",X"6C",X"63",
		X"FF",X"2A",X"A1",X"2F",X"11",X"B1",X"7F",X"2B",
		X"CC",X"59",X"30",X"F0",X"CC",X"11",X"AF",X"7F",
		X"2B",X"D6",X"11",X"5F",X"6D",X"2B",X"D8",X"75",
		X"CF",X"6C",X"63",X"11",X"B4",X"7F",X"2B",X"CC",
		X"59",X"31",X"F0",X"CC",X"11",X"B2",X"7F",X"2B",
		X"D6",X"11",X"3A",X"6D",X"2B",X"D8",X"75",X"CF",
		X"6C",X"63",X"FF",X"2B",X"A1",X"35",X"11",X"A2",
		X"7F",X"2B",X"CC",X"59",X"06",X"5E",X"9A",X"59",
		X"30",X"F0",X"CC",X"93",X"CC",X"1A",X"9A",X"E6",
		X"01",X"5E",X"9A",X"35",X"72",X"A8",X"11",X"A1",
		X"7F",X"2B",X"D6",X"11",X"44",X"6D",X"2B",X"D8",
		X"75",X"CF",X"6C",X"63",X"11",X"A8",X"7F",X"2B",
		X"D6",X"11",X"44",X"16",X"2B",X"D8",X"75",X"CF",
		X"6C",X"63",X"FF",X"2C",X"A1",X"1E",X"11",X"B1",
		X"7F",X"2B",X"CC",X"AD",X"E3",X"01",X"5E",X"9A",
		X"8C",X"3A",X"35",X"3F",X"BC",X"1A",X"9A",X"F0",
		X"CC",X"11",X"B4",X"7F",X"2B",X"CC",X"AD",X"E3",
		X"01",X"F0",X"CC",X"FF",X"2D",X"A1",X"2A",X"21",
		X"B0",X"2B",X"A4",X"00",X"FD",X"04",X"68",X"18",
		X"21",X"B2",X"2B",X"A6",X"21",X"B4",X"2B",X"AE",
		X"21",X"B6",X"2B",X"9C",X"21",X"B8",X"2B",X"9E",
		X"FF",X"21",X"A4",X"2B",X"B0",X"21",X"A6",X"2B",
		X"B2",X"21",X"AE",X"2B",X"B4",X"21",X"9C",X"2B",
		X"B6",X"21",X"9E",X"2B",X"B8",X"FF",X"2E",X"A1",
		X"3D",X"11",X"00",X"00",X"2B",X"3C",X"2B",X"40",
		X"2B",X"42",X"11",X"FC",X"01",X"2B",X"3E",X"2B",
		X"44",X"11",X"A1",X"35",X"2B",X"3A",X"59",X"04",
		X"5E",X"9A",X"59",X"FA",X"5E",X"44",X"11",X"00",
		X"02",X"F3",X"44",X"93",X"44",X"93",X"44",X"11",
		X"00",X"00",X"F3",X"44",X"93",X"44",X"93",X"44",
		X"F3",X"44",X"93",X"45",X"1A",X"9A",X"E6",X"01",
		X"5E",X"9A",X"35",X"72",X"B8",X"FF",X"2F",X"A1",
		X"42",X"59",X"05",X"5E",X"2C",X"1A",X"0E",X"B8",
		X"40",X"35",X"3F",X"AB",X"FF",X"75",X"21",X"3A",
		X"AD",X"2B",X"3C",X"21",X"3A",X"E3",X"01",X"2B",
		X"3A",X"59",X"F0",X"F8",X"3C",X"8C",X"90",X"35",
		X"72",X"C4",X"CF",X"68",X"90",X"AC",X"8C",X"10",
		X"35",X"72",X"CD",X"CF",X"66",X"90",X"AC",X"8C",
		X"50",X"35",X"72",X"D9",X"21",X"3A",X"F6",X"2B",
		X"3A",X"90",X"AC",X"1A",X"0E",X"99",X"3C",X"5E",
		X"40",X"63",X"FF",X"30",X"A1",X"4A",X"11",X"00",
		X"09",X"2B",X"44",X"21",X"3A",X"AD",X"E6",X"0B",
		X"E9",X"99",X"44",X"2B",X"44",X"7F",X"00",X"5E",
		X"42",X"21",X"44",X"7F",X"01",X"5E",X"43",X"21",
		X"3C",X"82",X"03",X"5E",X"45",X"59",X"00",X"5E",
		X"44",X"21",X"44",X"99",X"3E",X"2B",X"44",X"21",
		X"42",X"F3",X"44",X"21",X"3A",X"E3",X"01",X"2B",
		X"3A",X"FF",X"21",X"3C",X"82",X"03",X"5E",X"45",
		X"59",X"00",X"5E",X"44",X"21",X"44",X"99",X"3E",
		X"2B",X"44",X"11",X"00",X"00",X"F3",X"44",X"FF",
		X"34",X"A1",X"32",X"00",X"FD",X"04",X"68",X"18",
		X"90",X"53",X"91",X"47",X"07",X"90",X"52",X"91",
		X"46",X"07",X"90",X"53",X"91",X"47",X"07",X"90",
		X"52",X"91",X"46",X"07",X"90",X"53",X"91",X"47",
		X"07",X"90",X"54",X"91",X"48",X"07",X"90",X"53",
		X"91",X"47",X"07",X"90",X"52",X"91",X"46",X"07",
		X"90",X"53",X"91",X"47",X"1E",X"80",X"81",X"D0",
		X"A1",X"35",X"35",X"A1",X"5D",X"20",X"90",X"4A",
		X"91",X"3B",X"92",X"4D",X"0D",X"90",X"3A",X"91",
		X"4B",X"92",X"4E",X"0D",X"90",X"3B",X"91",X"4A",
		X"92",X"4D",X"0D",X"90",X"3A",X"91",X"4B",X"92",
		X"4E",X"0D",X"90",X"36",X"91",X"46",X"92",X"4B",
		X"0D",X"90",X"27",X"91",X"4E",X"92",X"57",X"0D",
		X"93",X"2A",X"80",X"81",X"82",X"0D",X"93",X"25",
		X"0D",X"90",X"4A",X"91",X"3B",X"92",X"4D",X"83",
		X"0D",X"90",X"3A",X"91",X"4B",X"92",X"4E",X"0D",
		X"90",X"3B",X"91",X"4A",X"92",X"4D",X"0D",X"90",
		X"3A",X"91",X"4B",X"92",X"4E",X"0D",X"90",X"36",
		X"91",X"46",X"92",X"4B",X"0D",X"90",X"27",X"D0",
		X"A1",X"36",X"36",X"A1",X"5A",X"91",X"4E",X"92",
		X"57",X"0D",X"93",X"2A",X"80",X"81",X"82",X"0D",
		X"93",X"25",X"0D",X"90",X"2E",X"83",X"0D",X"91",
		X"4A",X"90",X"53",X"92",X"35",X"0D",X"90",X"2E",
		X"81",X"82",X"0D",X"91",X"4A",X"90",X"52",X"92",
		X"29",X"0D",X"90",X"29",X"81",X"82",X"0D",X"91",
		X"48",X"90",X"50",X"92",X"29",X"0D",X"90",X"29",
		X"81",X"82",X"0D",X"91",X"48",X"90",X"50",X"92",
		X"35",X"0D",X"90",X"48",X"91",X"2C",X"92",X"50",
		X"06",X"90",X"4A",X"92",X"52",X"06",X"90",X"36",
		X"91",X"48",X"92",X"50",X"0D",X"90",X"2C",X"91",
		X"48",X"92",X"50",X"0D",X"D0",X"A1",X"37",X"37",
		X"A1",X"5B",X"90",X"36",X"91",X"47",X"92",X"4B",
		X"0D",X"90",X"2E",X"00",X"FD",X"04",X"68",X"18",
		X"91",X"4A",X"92",X"4D",X"0D",X"80",X"81",X"82",
		X"26",X"90",X"3B",X"91",X"4B",X"92",X"4E",X"0D",
		X"90",X"3A",X"91",X"4D",X"92",X"50",X"0D",X"90",
		X"3B",X"91",X"4B",X"92",X"4E",X"0D",X"90",X"3A",
		X"91",X"4D",X"92",X"50",X"0D",X"90",X"2E",X"91",
		X"4A",X"92",X"4D",X"0D",X"90",X"2E",X"91",X"56",
		X"92",X"59",X"0D",X"93",X"2A",X"80",X"81",X"82",
		X"0D",X"93",X"25",X"0D",X"90",X"4B",X"91",X"3B",
		X"92",X"4E",X"83",X"0D",X"90",X"3A",X"91",X"4D",
		X"92",X"50",X"0D",X"90",X"3B",X"91",X"4B",X"D0",
		X"A1",X"38",X"38",X"A1",X"5A",X"92",X"4E",X"0D",
		X"90",X"3A",X"91",X"4D",X"92",X"50",X"0D",X"90",
		X"2E",X"91",X"4A",X"92",X"4D",X"0D",X"90",X"2E",
		X"91",X"56",X"92",X"59",X"0D",X"93",X"2A",X"80",
		X"81",X"82",X"0D",X"93",X"25",X"0D",X"90",X"2C",
		X"83",X"0D",X"91",X"57",X"90",X"5A",X"92",X"35",
		X"0D",X"90",X"2C",X"81",X"82",X"0D",X"91",X"56",
		X"90",X"59",X"92",X"35",X"0D",X"90",X"2E",X"81",
		X"82",X"0D",X"91",X"52",X"90",X"57",X"92",X"36",
		X"0D",X"90",X"2E",X"81",X"82",X"0D",X"91",X"52",
		X"90",X"57",X"92",X"36",X"0D",X"90",X"2F",X"81",
		X"82",X"0D",X"91",X"53",X"D0",X"A1",X"39",X"39",
		X"A1",X"5A",X"90",X"57",X"92",X"38",X"06",X"90",
		X"56",X"91",X"59",X"06",X"90",X"2F",X"91",X"53",
		X"92",X"57",X"06",X"81",X"82",X"06",X"90",X"52",
		X"91",X"38",X"92",X"56",X"06",X"80",X"82",X"06",
		X"90",X"4F",X"91",X"33",X"92",X"57",X"06",X"80",
		X"82",X"06",X"81",X"26",X"90",X"43",X"91",X"33",
		X"92",X"46",X"06",X"90",X"44",X"92",X"48",X"06",
		X"93",X"25",X"90",X"33",X"91",X"43",X"92",X"46",
		X"0D",X"80",X"83",X"0D",X"90",X"33",X"93",X"2C",
		X"81",X"82",X"0D",X"00",X"FD",X"04",X"68",X"18",
		X"90",X"33",X"93",X"2C",X"0D",X"90",X"33",X"93",
		X"25",X"0D",X"91",X"43",X"90",X"4B",X"D0",X"A1",
		X"3A",X"3A",X"A1",X"59",X"83",X"0D",X"92",X"33",
		X"93",X"2C",X"0D",X"90",X"44",X"91",X"33",X"93",
		X"2C",X"92",X"48",X"0D",X"91",X"33",X"93",X"25",
		X"0D",X"80",X"81",X"82",X"83",X"0D",X"90",X"33",
		X"93",X"2C",X"0D",X"90",X"33",X"93",X"2C",X"0D",
		X"90",X"33",X"93",X"25",X"0D",X"80",X"83",X"0D",
		X"90",X"33",X"93",X"2C",X"0D",X"91",X"41",X"90",
		X"44",X"92",X"2E",X"93",X"2C",X"06",X"90",X"43",
		X"91",X"46",X"06",X"90",X"2E",X"93",X"25",X"91",
		X"41",X"92",X"44",X"0D",X"80",X"83",X"0D",X"90",
		X"2E",X"93",X"2C",X"81",X"82",X"0D",X"90",X"2E",
		X"93",X"2C",X"D0",X"A1",X"3B",X"3B",X"A1",X"5A",
		X"0D",X"90",X"2E",X"93",X"25",X"0D",X"91",X"41",
		X"90",X"4A",X"83",X"0D",X"92",X"2E",X"93",X"2C",
		X"0D",X"90",X"43",X"91",X"33",X"93",X"2C",X"92",
		X"4A",X"06",X"92",X"4B",X"06",X"91",X"33",X"93",
		X"25",X"92",X"46",X"0D",X"80",X"81",X"83",X"0D",
		X"90",X"33",X"93",X"2C",X"82",X"0D",X"90",X"33",
		X"93",X"2C",X"0D",X"90",X"33",X"93",X"25",X"0D",
		X"80",X"83",X"0D",X"90",X"33",X"93",X"2C",X"0D",
		X"91",X"3F",X"90",X"43",X"92",X"33",X"93",X"2C",
		X"06",X"90",X"3C",X"91",X"46",X"06",X"90",X"33",
		X"93",X"25",X"91",X"3A",X"92",X"43",X"0D",X"D0",
		X"A1",X"3C",X"3C",X"A1",X"5B",X"80",X"83",X"0D",
		X"90",X"33",X"93",X"2C",X"81",X"82",X"0D",X"90",
		X"33",X"93",X"2C",X"0D",X"90",X"33",X"93",X"25",
		X"0D",X"91",X"43",X"90",X"46",X"83",X"0D",X"92",
		X"33",X"93",X"2C",X"0D",X"90",X"3E",X"91",X"2C",
		X"93",X"2C",X"92",X"46",X"06",X"90",X"3F",X"92",
		X"48",X"06",X"90",X"00",X"FD",X"04",X"68",X"18",
		X"2C",X"93",X"25",X"91",X"3C",X"92",X"44",X"0D",
		X"80",X"83",X"0D",X"90",X"2C",X"93",X"2C",X"81",
		X"82",X"0D",X"90",X"2C",X"93",X"2C",X"0D",X"90",
		X"2C",X"93",X"25",X"0D",X"80",X"83",X"0D",X"90",
		X"2C",X"93",X"2C",X"0D",X"91",X"3A",X"90",X"3E",
		X"92",X"2E",X"D0",X"A1",X"3D",X"3D",X"A1",X"59",
		X"93",X"2C",X"06",X"90",X"3C",X"91",X"3F",X"06",
		X"90",X"2E",X"93",X"25",X"91",X"3A",X"92",X"3E",
		X"0D",X"80",X"83",X"0D",X"90",X"2E",X"93",X"2C",
		X"81",X"82",X"0D",X"90",X"2E",X"93",X"2C",X"0D",
		X"90",X"2E",X"93",X"25",X"0D",X"91",X"38",X"90",
		X"41",X"83",X"0D",X"92",X"2E",X"93",X"2C",X"0D",
		X"90",X"3B",X"91",X"33",X"93",X"2C",X"92",X"44",
		X"0D",X"91",X"33",X"93",X"25",X"0D",X"80",X"81",
		X"82",X"83",X"0D",X"90",X"3A",X"91",X"33",X"93",
		X"2C",X"92",X"43",X"0D",X"91",X"33",X"93",X"2C",
		X"0D",X"90",X"33",X"93",X"25",X"81",X"D0",X"A1",
		X"3E",X"3E",X"A1",X"5B",X"82",X"0D",X"80",X"83",
		X"0D",X"90",X"33",X"93",X"2C",X"0D",X"91",X"4F",
		X"90",X"46",X"92",X"33",X"93",X"2C",X"06",X"90",
		X"48",X"06",X"90",X"33",X"93",X"25",X"92",X"46",
		X"0D",X"80",X"83",X"0D",X"90",X"33",X"93",X"2C",
		X"91",X"50",X"82",X"0D",X"90",X"33",X"93",X"2C",
		X"0D",X"90",X"33",X"93",X"25",X"0D",X"90",X"4F",
		X"91",X"4B",X"83",X"0D",X"92",X"33",X"93",X"2C",
		X"0D",X"90",X"52",X"91",X"2C",X"93",X"2C",X"92",
		X"48",X"0D",X"91",X"2C",X"93",X"25",X"0D",X"81",
		X"82",X"83",X"0D",X"90",X"2C",X"93",X"2C",X"91",
		X"50",X"0D",X"90",X"2C",X"D0",X"A1",X"3F",X"3F",
		X"A1",X"59",X"93",X"2C",X"0D",X"90",X"2C",X"93",
		X"25",X"81",X"0D",X"80",X"83",X"0D",X"90",X"2C",
		X"93",X"2C",X"0D",X"00",X"FD",X"04",X"68",X"18",
		X"91",X"4B",X"90",X"44",X"92",X"2E",X"93",X"2C",
		X"06",X"90",X"46",X"06",X"90",X"2E",X"93",X"25",
		X"92",X"44",X"0D",X"80",X"83",X"0D",X"90",X"2E",
		X"93",X"2C",X"91",X"4D",X"82",X"0D",X"90",X"2E",
		X"93",X"2C",X"0D",X"90",X"2E",X"93",X"25",X"0D",
		X"90",X"4F",X"91",X"4A",X"83",X"0D",X"92",X"2E",
		X"93",X"2C",X"0D",X"90",X"50",X"91",X"33",X"93",
		X"2C",X"92",X"4A",X"06",X"92",X"4B",X"06",X"91",
		X"33",X"93",X"25",X"92",X"46",X"D0",X"A1",X"40",
		X"40",X"A1",X"5A",X"0D",X"81",X"83",X"0D",X"90",
		X"33",X"93",X"2C",X"91",X"4F",X"82",X"0D",X"90",
		X"32",X"93",X"2C",X"0D",X"90",X"32",X"93",X"25",
		X"81",X"0D",X"80",X"83",X"0D",X"90",X"32",X"93",
		X"2C",X"0D",X"91",X"4B",X"90",X"43",X"92",X"30",
		X"93",X"2C",X"06",X"90",X"46",X"06",X"90",X"30",
		X"93",X"25",X"92",X"43",X"0D",X"80",X"83",X"0D",
		X"90",X"30",X"93",X"2C",X"91",X"4A",X"82",X"0D",
		X"90",X"2E",X"93",X"2C",X"0D",X"90",X"4A",X"91",
		X"2E",X"93",X"25",X"0D",X"92",X"46",X"81",X"83",
		X"0D",X"91",X"2E",X"93",X"2C",X"0D",X"90",X"4F",
		X"91",X"2C",X"D0",X"A1",X"41",X"41",X"A1",X"5A",
		X"93",X"2C",X"92",X"46",X"06",X"92",X"48",X"06",
		X"91",X"2C",X"93",X"25",X"92",X"44",X"0D",X"81",
		X"83",X"0D",X"90",X"2C",X"93",X"2C",X"91",X"4D",
		X"82",X"0D",X"90",X"2C",X"93",X"2C",X"0D",X"90",
		X"2C",X"93",X"25",X"81",X"0D",X"91",X"48",X"80",
		X"83",X"0D",X"90",X"2C",X"93",X"2C",X"0D",X"90",
		X"50",X"91",X"2E",X"93",X"2C",X"92",X"3E",X"06",
		X"92",X"3F",X"06",X"91",X"2E",X"93",X"25",X"92",
		X"3E",X"0D",X"81",X"83",X"0D",X"90",X"2E",X"93",
		X"2C",X"91",X"52",X"82",X"0D",X"90",X"2E",X"93",
		X"2C",X"0D",X"90",X"00",X"FD",X"04",X"68",X"18",
		X"2E",X"93",X"25",X"0D",X"D0",X"A1",X"42",X"42",
		X"A1",X"3D",X"90",X"50",X"91",X"41",X"83",X"0D",
		X"92",X"2E",X"93",X"2C",X"0D",X"91",X"4D",X"92",
		X"33",X"93",X"2C",X"0D",X"90",X"33",X"93",X"25",
		X"82",X"0D",X"80",X"83",X"0D",X"90",X"33",X"93",
		X"2C",X"91",X"4B",X"92",X"43",X"0D",X"90",X"33",
		X"93",X"2C",X"0D",X"90",X"33",X"93",X"25",X"81",
		X"82",X"0D",X"80",X"83",X"0D",X"90",X"33",X"93",
		X"25",X"0D",X"80",X"83",X"D0",X"A1",X"43",X"43",
		X"A1",X"5D",X"90",X"47",X"91",X"28",X"92",X"4C",
		X"0C",X"93",X"20",X"91",X"34",X"0C",X"90",X"44",
		X"91",X"28",X"92",X"47",X"83",X"0C",X"93",X"20",
		X"91",X"34",X"90",X"45",X"92",X"48",X"0C",X"91",
		X"28",X"90",X"47",X"92",X"4A",X"83",X"0C",X"93",
		X"20",X"91",X"34",X"06",X"93",X"20",X"06",X"90",
		X"45",X"91",X"28",X"92",X"48",X"83",X"0C",X"93",
		X"20",X"91",X"34",X"90",X"44",X"92",X"47",X"06",
		X"83",X"06",X"90",X"40",X"91",X"2D",X"92",X"45",
		X"0C",X"93",X"20",X"91",X"39",X"0C",X"90",X"40",
		X"91",X"2D",X"92",X"45",X"83",X"0C",X"93",X"20",
		X"91",X"39",X"90",X"45",X"D0",X"A1",X"44",X"44",
		X"A1",X"5B",X"92",X"48",X"0C",X"91",X"2D",X"90",
		X"48",X"92",X"4C",X"83",X"0C",X"93",X"20",X"91",
		X"39",X"0C",X"90",X"20",X"92",X"47",X"91",X"2D",
		X"93",X"4A",X"06",X"80",X"06",X"90",X"20",X"92",
		X"45",X"91",X"39",X"93",X"48",X"0C",X"91",X"2C",
		X"90",X"44",X"92",X"47",X"83",X"0C",X"93",X"20",
		X"91",X"38",X"0C",X"91",X"2C",X"83",X"0C",X"93",
		X"20",X"90",X"45",X"91",X"38",X"92",X"48",X"0C",
		X"91",X"28",X"90",X"47",X"92",X"4A",X"83",X"0C",
		X"93",X"20",X"91",X"34",X"06",X"93",X"20",X"06",
		X"90",X"47",X"91",X"00",X"FD",X"04",X"68",X"18",
		X"28",X"92",X"4C",X"83",X"0C",X"93",X"20",X"D0",
		X"A1",X"45",X"45",X"A1",X"59",X"91",X"34",X"06",
		X"83",X"06",X"90",X"45",X"91",X"2D",X"92",X"48",
		X"0C",X"93",X"20",X"91",X"39",X"0C",X"90",X"40",
		X"91",X"2D",X"92",X"45",X"83",X"0C",X"93",X"20",
		X"91",X"39",X"0C",X"90",X"40",X"91",X"2D",X"92",
		X"45",X"83",X"0C",X"93",X"20",X"91",X"39",X"0C",
		X"90",X"20",X"91",X"2F",X"82",X"83",X"06",X"80",
		X"06",X"90",X"20",X"91",X"30",X"0C",X"91",X"32",
		X"80",X"0C",X"90",X"20",X"92",X"41",X"93",X"4A",
		X"91",X"26",X"0C",X"80",X"81",X"82",X"83",X"0C",
		X"90",X"20",X"92",X"45",X"91",X"26",X"93",X"4D",
		X"0C",X"90",X"48",X"D0",X"A1",X"46",X"46",X"A1",
		X"5A",X"92",X"51",X"81",X"83",X"0C",X"91",X"26",
		X"93",X"20",X"90",X"48",X"06",X"91",X"26",X"90",
		X"20",X"93",X"48",X"06",X"91",X"2D",X"90",X"47",
		X"92",X"4F",X"83",X"0C",X"93",X"20",X"91",X"29",
		X"90",X"45",X"92",X"4D",X"06",X"83",X"06",X"90",
		X"43",X"91",X"24",X"92",X"4C",X"0C",X"93",X"20",
		X"91",X"30",X"80",X"82",X"0C",X"81",X"83",X"0C",
		X"90",X"20",X"92",X"40",X"91",X"30",X"93",X"48",
		X"0C",X"90",X"43",X"92",X"4C",X"81",X"83",X"0C",
		X"91",X"24",X"93",X"20",X"90",X"45",X"06",X"91",
		X"25",X"90",X"43",X"06",X"91",X"26",X"90",X"20",
		X"D0",X"A1",X"47",X"47",X"A1",X"5B",X"92",X"41",
		X"93",X"4A",X"06",X"80",X"06",X"90",X"20",X"92",
		X"40",X"91",X"27",X"93",X"48",X"0C",X"90",X"44",
		X"92",X"47",X"81",X"83",X"0C",X"91",X"3B",X"93",
		X"20",X"80",X"0C",X"90",X"44",X"92",X"47",X"81",
		X"83",X"0C",X"91",X"3B",X"93",X"20",X"90",X"45",
		X"92",X"48",X"0C",X"90",X"47",X"92",X"4A",X"81",
		X"83",X"0C",X"91",X"00",X"FD",X"04",X"68",X"18",
		X"34",X"93",X"20",X"06",X"93",X"20",X"06",X"90",
		X"47",X"92",X"4C",X"81",X"83",X"0C",X"91",X"38",
		X"93",X"20",X"06",X"83",X"06",X"90",X"45",X"91",
		X"2D",X"92",X"48",X"0C",X"93",X"20",X"91",X"34",
		X"0C",X"90",X"40",X"D0",X"A1",X"48",X"48",X"A1",
		X"59",X"91",X"2D",X"92",X"45",X"83",X"0C",X"93",
		X"20",X"91",X"34",X"0C",X"90",X"40",X"91",X"2D",
		X"92",X"45",X"83",X"0C",X"93",X"20",X"81",X"0C",
		X"90",X"20",X"82",X"83",X"06",X"80",X"06",X"90",
		X"20",X"0C",X"92",X"47",X"91",X"28",X"90",X"4C",
		X"0C",X"93",X"20",X"91",X"34",X"0C",X"90",X"44",
		X"91",X"28",X"92",X"47",X"83",X"0C",X"93",X"20",
		X"91",X"34",X"90",X"45",X"92",X"48",X"0C",X"91",
		X"28",X"90",X"47",X"92",X"4A",X"83",X"0C",X"93",
		X"20",X"91",X"34",X"06",X"93",X"20",X"06",X"90",
		X"45",X"91",X"28",X"92",X"48",X"83",X"0C",X"D0",
		X"A1",X"49",X"49",X"A1",X"5B",X"93",X"20",X"91",
		X"34",X"90",X"44",X"92",X"47",X"06",X"83",X"06",
		X"90",X"40",X"91",X"2D",X"92",X"45",X"0C",X"93",
		X"20",X"91",X"39",X"0C",X"90",X"40",X"91",X"2D",
		X"92",X"45",X"83",X"0C",X"93",X"20",X"91",X"39",
		X"90",X"45",X"92",X"48",X"0C",X"91",X"2D",X"90",
		X"48",X"92",X"4C",X"83",X"0C",X"93",X"20",X"91",
		X"39",X"0C",X"90",X"20",X"92",X"47",X"91",X"2D",
		X"93",X"4A",X"06",X"80",X"06",X"90",X"20",X"92",
		X"45",X"91",X"39",X"93",X"48",X"0C",X"91",X"2C",
		X"90",X"44",X"92",X"47",X"83",X"0C",X"93",X"20",
		X"91",X"38",X"0C",X"91",X"2C",X"D0",X"A1",X"4A",
		X"4A",X"A1",X"59",X"83",X"0C",X"93",X"20",X"90",
		X"45",X"91",X"38",X"92",X"48",X"0C",X"91",X"28",
		X"90",X"47",X"92",X"4A",X"83",X"0C",X"93",X"20",
		X"91",X"34",X"06",X"00",X"FD",X"04",X"68",X"18",
		X"93",X"20",X"06",X"90",X"47",X"91",X"28",X"92",
		X"4C",X"83",X"0C",X"93",X"20",X"91",X"34",X"06",
		X"83",X"06",X"90",X"45",X"91",X"2D",X"92",X"48",
		X"0C",X"93",X"20",X"91",X"39",X"0C",X"90",X"40",
		X"91",X"2D",X"92",X"45",X"83",X"0C",X"93",X"20",
		X"91",X"39",X"0C",X"90",X"40",X"91",X"2D",X"92",
		X"45",X"83",X"0C",X"93",X"20",X"91",X"39",X"0C",
		X"90",X"20",X"91",X"2F",X"82",X"83",X"D0",X"A1",
		X"4B",X"4B",X"A1",X"5A",X"06",X"80",X"06",X"90",
		X"20",X"91",X"30",X"0C",X"91",X"32",X"80",X"0C",
		X"90",X"20",X"92",X"41",X"93",X"4A",X"91",X"26",
		X"0C",X"80",X"81",X"82",X"83",X"0C",X"90",X"20",
		X"92",X"45",X"91",X"26",X"93",X"4D",X"0C",X"90",
		X"48",X"92",X"51",X"81",X"83",X"0C",X"91",X"26",
		X"93",X"20",X"90",X"48",X"06",X"91",X"26",X"90",
		X"20",X"93",X"48",X"06",X"91",X"2D",X"90",X"47",
		X"92",X"4F",X"83",X"0C",X"93",X"20",X"91",X"29",
		X"90",X"45",X"92",X"4D",X"06",X"83",X"06",X"90",
		X"43",X"91",X"24",X"92",X"4C",X"0C",X"93",X"20",
		X"91",X"30",X"80",X"D0",X"A1",X"4C",X"4C",X"A1",
		X"5A",X"82",X"0C",X"81",X"83",X"0C",X"90",X"20",
		X"92",X"40",X"91",X"30",X"93",X"48",X"0C",X"90",
		X"43",X"92",X"4C",X"81",X"83",X"0C",X"91",X"24",
		X"93",X"20",X"90",X"45",X"06",X"91",X"25",X"90",
		X"43",X"06",X"91",X"26",X"90",X"20",X"92",X"41",
		X"93",X"4A",X"06",X"80",X"06",X"90",X"20",X"92",
		X"40",X"91",X"27",X"93",X"48",X"0C",X"90",X"44",
		X"92",X"47",X"81",X"83",X"0C",X"91",X"3B",X"93",
		X"20",X"80",X"0C",X"90",X"44",X"92",X"47",X"81",
		X"83",X"0C",X"91",X"3B",X"93",X"20",X"90",X"45",
		X"92",X"48",X"0C",X"90",X"47",X"92",X"4A",X"81",
		X"D0",X"A1",X"4D",X"00",X"FD",X"04",X"68",X"18",
		X"4D",X"A1",X"5A",X"83",X"0C",X"91",X"34",X"93",
		X"20",X"06",X"93",X"20",X"06",X"90",X"47",X"92",
		X"4C",X"81",X"83",X"0C",X"91",X"38",X"93",X"20",
		X"06",X"83",X"06",X"90",X"45",X"91",X"2D",X"92",
		X"48",X"0C",X"93",X"20",X"91",X"34",X"0C",X"90",
		X"40",X"91",X"2D",X"92",X"45",X"83",X"0C",X"93",
		X"20",X"91",X"34",X"0C",X"90",X"40",X"91",X"2D",
		X"92",X"45",X"83",X"0C",X"93",X"20",X"81",X"0C",
		X"90",X"20",X"82",X"83",X"06",X"80",X"06",X"90",
		X"20",X"0C",X"91",X"39",X"92",X"45",X"90",X"40",
		X"0C",X"92",X"20",X"93",X"4C",X"0C",X"92",X"45",
		X"83",X"0C",X"D0",X"A1",X"4E",X"4E",X"A1",X"5A",
		X"93",X"20",X"92",X"4C",X"0C",X"90",X"3C",X"92",
		X"45",X"83",X"0C",X"93",X"20",X"92",X"4C",X"06",
		X"93",X"20",X"06",X"92",X"45",X"83",X"0C",X"93",
		X"20",X"92",X"4C",X"06",X"83",X"06",X"90",X"38",
		X"92",X"44",X"91",X"3E",X"0C",X"92",X"20",X"93",
		X"4C",X"0C",X"92",X"44",X"83",X"0C",X"93",X"20",
		X"92",X"4C",X"0C",X"91",X"3B",X"92",X"44",X"83",
		X"0C",X"93",X"20",X"92",X"4C",X"0C",X"92",X"20",
		X"93",X"44",X"06",X"82",X"06",X"92",X"20",X"93",
		X"4C",X"0C",X"90",X"39",X"92",X"45",X"91",X"3C",
		X"83",X"0C",X"92",X"20",X"93",X"4C",X"0C",X"D0",
		X"A1",X"4F",X"4F",X"A1",X"5B",X"92",X"45",X"83",
		X"0C",X"93",X"20",X"92",X"4C",X"0C",X"90",X"34",
		X"92",X"45",X"91",X"39",X"83",X"0C",X"92",X"20",
		X"93",X"4C",X"06",X"92",X"20",X"06",X"92",X"45",
		X"83",X"0C",X"93",X"20",X"92",X"4C",X"06",X"83",
		X"06",X"91",X"38",X"92",X"44",X"0C",X"93",X"20",
		X"92",X"4C",X"0C",X"92",X"44",X"83",X"0C",X"93",
		X"20",X"92",X"4C",X"0C",X"90",X"3B",X"92",X"44",
		X"83",X"0C",X"93",X"00",X"FD",X"04",X"68",X"18",
		X"20",X"92",X"4C",X"0C",X"92",X"20",X"93",X"44",
		X"06",X"82",X"06",X"92",X"20",X"93",X"4C",X"0C",
		X"90",X"39",X"92",X"45",X"91",X"40",X"83",X"0C",
		X"92",X"20",X"D0",X"A1",X"50",X"50",X"A1",X"5A",
		X"93",X"4C",X"0C",X"92",X"45",X"83",X"0C",X"93",
		X"20",X"92",X"4C",X"0C",X"91",X"3C",X"92",X"45",
		X"83",X"0C",X"93",X"20",X"92",X"4C",X"06",X"93",
		X"20",X"06",X"92",X"45",X"83",X"0C",X"93",X"20",
		X"92",X"4C",X"06",X"83",X"06",X"90",X"38",X"92",
		X"44",X"91",X"3E",X"0C",X"92",X"20",X"93",X"4C",
		X"0C",X"92",X"44",X"83",X"0C",X"93",X"20",X"92",
		X"4C",X"0C",X"91",X"3B",X"92",X"44",X"83",X"0C",
		X"93",X"20",X"92",X"4C",X"0C",X"92",X"20",X"93",
		X"44",X"06",X"82",X"06",X"92",X"20",X"93",X"4C",
		X"0C",X"90",X"39",X"92",X"45",X"91",X"3C",X"D0",
		X"A1",X"51",X"51",X"A1",X"59",X"83",X"0C",X"92",
		X"20",X"93",X"4C",X"0C",X"91",X"40",X"92",X"45",
		X"83",X"0C",X"93",X"20",X"92",X"4C",X"0C",X"91",
		X"45",X"92",X"45",X"83",X"0C",X"93",X"20",X"92",
		X"4C",X"06",X"93",X"20",X"06",X"91",X"45",X"92",
		X"45",X"83",X"0C",X"93",X"20",X"92",X"4C",X"06",
		X"83",X"06",X"90",X"3E",X"92",X"44",X"91",X"44",
		X"0C",X"92",X"20",X"93",X"4C",X"0C",X"92",X"44",
		X"83",X"0C",X"93",X"20",X"92",X"4C",X"0C",X"92",
		X"44",X"83",X"0C",X"93",X"20",X"92",X"4C",X"0C",
		X"92",X"20",X"93",X"44",X"06",X"82",X"06",X"92",
		X"20",X"93",X"4C",X"D0",X"A1",X"52",X"52",X"A1",
		X"5A",X"0C",X"92",X"47",X"93",X"4C",X"80",X"81",
		X"0C",X"90",X"20",X"91",X"34",X"0C",X"90",X"47",
		X"91",X"28",X"92",X"44",X"83",X"0C",X"93",X"20",
		X"91",X"34",X"90",X"45",X"92",X"48",X"0C",X"91",
		X"28",X"90",X"47",X"00",X"FD",X"04",X"68",X"18",
		X"92",X"4A",X"83",X"0C",X"93",X"20",X"91",X"34",
		X"06",X"93",X"20",X"06",X"90",X"48",X"91",X"28",
		X"92",X"45",X"83",X"0C",X"93",X"20",X"91",X"34",
		X"90",X"44",X"92",X"47",X"06",X"83",X"06",X"90",
		X"40",X"91",X"2D",X"92",X"45",X"0C",X"93",X"20",
		X"91",X"39",X"0C",X"90",X"40",X"91",X"2D",X"92",
		X"45",X"83",X"0C",X"93",X"20",X"D0",X"A1",X"53",
		X"53",X"A1",X"5B",X"91",X"39",X"90",X"48",X"92",
		X"45",X"0C",X"91",X"2D",X"90",X"4C",X"92",X"48",
		X"83",X"0C",X"93",X"20",X"91",X"39",X"0C",X"90",
		X"20",X"92",X"47",X"91",X"2D",X"93",X"4A",X"06",
		X"80",X"06",X"90",X"20",X"92",X"45",X"91",X"39",
		X"93",X"48",X"0C",X"91",X"2C",X"90",X"44",X"92",
		X"47",X"83",X"0C",X"93",X"20",X"91",X"38",X"0C",
		X"91",X"2C",X"83",X"0C",X"93",X"20",X"90",X"48",
		X"91",X"38",X"92",X"45",X"0C",X"91",X"28",X"90",
		X"47",X"92",X"4A",X"83",X"0C",X"93",X"20",X"91",
		X"34",X"06",X"93",X"20",X"06",X"90",X"4C",X"91",
		X"28",X"92",X"47",X"D0",X"A1",X"54",X"54",X"A1",
		X"5A",X"83",X"0C",X"93",X"20",X"91",X"34",X"06",
		X"83",X"06",X"90",X"45",X"91",X"2D",X"92",X"48",
		X"0C",X"93",X"20",X"91",X"39",X"0C",X"90",X"40",
		X"91",X"2D",X"92",X"45",X"83",X"0C",X"93",X"20",
		X"91",X"39",X"0C",X"90",X"40",X"91",X"2D",X"92",
		X"45",X"83",X"0C",X"93",X"20",X"91",X"39",X"0C",
		X"90",X"20",X"91",X"2F",X"82",X"83",X"06",X"80",
		X"06",X"90",X"20",X"91",X"30",X"0C",X"91",X"32",
		X"80",X"0C",X"90",X"20",X"92",X"4A",X"93",X"41",
		X"91",X"26",X"0C",X"80",X"81",X"82",X"83",X"0C",
		X"90",X"20",X"92",X"45",X"91",X"26",X"93",X"4D",
		X"D0",X"A1",X"55",X"55",X"A1",X"59",X"0C",X"90",
		X"48",X"92",X"51",X"00",X"FD",X"04",X"68",X"18",
		X"81",X"83",X"0C",X"91",X"26",X"93",X"20",X"90",
		X"48",X"06",X"91",X"26",X"90",X"20",X"93",X"48",
		X"06",X"91",X"2D",X"90",X"4F",X"92",X"47",X"83",
		X"0C",X"93",X"20",X"91",X"29",X"90",X"4D",X"92",
		X"45",X"06",X"83",X"06",X"90",X"43",X"91",X"24",
		X"92",X"4C",X"0C",X"93",X"20",X"91",X"30",X"80",
		X"82",X"0C",X"81",X"83",X"0C",X"90",X"20",X"92",
		X"40",X"91",X"30",X"93",X"48",X"0C",X"90",X"4C",
		X"92",X"43",X"81",X"83",X"0C",X"91",X"24",X"93",
		X"20",X"92",X"45",X"06",X"91",X"25",X"92",X"43",
		X"06",X"D0",X"A1",X"56",X"56",X"A1",X"5A",X"91",
		X"26",X"90",X"20",X"92",X"41",X"93",X"4A",X"06",
		X"80",X"06",X"90",X"20",X"92",X"48",X"91",X"27",
		X"93",X"40",X"0C",X"90",X"44",X"92",X"47",X"81",
		X"83",X"0C",X"91",X"3B",X"93",X"20",X"80",X"0C",
		X"90",X"44",X"92",X"47",X"81",X"83",X"0C",X"91",
		X"3B",X"93",X"20",X"90",X"48",X"92",X"45",X"0C",
		X"90",X"47",X"92",X"4A",X"81",X"83",X"0C",X"91",
		X"34",X"93",X"20",X"06",X"93",X"20",X"06",X"90",
		X"47",X"92",X"4C",X"81",X"83",X"0C",X"91",X"38",
		X"93",X"20",X"06",X"83",X"06",X"90",X"45",X"91",
		X"2D",X"92",X"48",X"0C",X"93",X"20",X"D0",X"A1",
		X"57",X"57",X"A1",X"5A",X"91",X"34",X"0C",X"90",
		X"45",X"91",X"2D",X"92",X"40",X"83",X"0C",X"93",
		X"20",X"91",X"34",X"0C",X"90",X"45",X"91",X"2D",
		X"92",X"40",X"83",X"0C",X"93",X"20",X"81",X"0C",
		X"90",X"20",X"82",X"83",X"06",X"80",X"06",X"90",
		X"20",X"0C",X"92",X"47",X"91",X"28",X"90",X"4C",
		X"0C",X"93",X"20",X"91",X"34",X"0C",X"90",X"44",
		X"91",X"28",X"92",X"47",X"83",X"0C",X"93",X"20",
		X"91",X"34",X"90",X"45",X"92",X"48",X"0C",X"91",
		X"28",X"90",X"4A",X"00",X"FD",X"04",X"68",X"18",
		X"92",X"47",X"83",X"0C",X"93",X"20",X"91",X"34",
		X"06",X"93",X"20",X"06",X"90",X"45",X"91",X"28",
		X"D0",X"A1",X"58",X"58",X"A1",X"5A",X"92",X"48",
		X"83",X"0C",X"93",X"20",X"91",X"34",X"90",X"47",
		X"92",X"44",X"06",X"83",X"06",X"90",X"40",X"91",
		X"2D",X"92",X"45",X"0C",X"93",X"20",X"91",X"39",
		X"0C",X"90",X"40",X"91",X"2D",X"92",X"45",X"83",
		X"0C",X"93",X"20",X"91",X"39",X"90",X"45",X"92",
		X"48",X"0C",X"91",X"2D",X"90",X"4C",X"92",X"48",
		X"83",X"0C",X"93",X"20",X"91",X"39",X"0C",X"90",
		X"20",X"92",X"4A",X"91",X"2D",X"93",X"47",X"06",
		X"80",X"06",X"90",X"20",X"92",X"45",X"91",X"39",
		X"93",X"48",X"0C",X"91",X"2C",X"90",X"47",X"92",
		X"44",X"83",X"0C",X"93",X"20",X"D0",X"A1",X"59",
		X"59",X"A1",X"5A",X"91",X"38",X"0C",X"91",X"2C",
		X"83",X"0C",X"93",X"20",X"90",X"45",X"91",X"38",
		X"92",X"48",X"0C",X"91",X"28",X"90",X"47",X"92",
		X"4A",X"83",X"0C",X"93",X"20",X"91",X"34",X"06",
		X"93",X"20",X"06",X"90",X"47",X"91",X"28",X"92",
		X"4C",X"83",X"0C",X"93",X"20",X"91",X"34",X"06",
		X"83",X"06",X"90",X"45",X"91",X"2D",X"92",X"48",
		X"0C",X"93",X"20",X"91",X"39",X"0C",X"90",X"40",
		X"91",X"2D",X"92",X"45",X"83",X"0C",X"93",X"20",
		X"91",X"39",X"0C",X"90",X"45",X"91",X"2D",X"92",
		X"40",X"83",X"0C",X"93",X"20",X"91",X"39",X"0C",
		X"90",X"20",X"D0",X"A1",X"5A",X"5A",X"A1",X"11",
		X"91",X"2F",X"82",X"83",X"06",X"80",X"06",X"90",
		X"20",X"91",X"30",X"0C",X"80",X"81",X"D0",X"A1",
		X"5B",X"5B",X"A1",X"5D",X"90",X"30",X"0B",X"91",
		X"3C",X"0B",X"91",X"3F",X"0B",X"91",X"43",X"0B",
		X"91",X"3F",X"80",X"0B",X"90",X"3C",X"81",X"0B",
		X"90",X"3F",X"0B",X"00",X"FD",X"04",X"68",X"18",
		X"90",X"3C",X"0B",X"90",X"37",X"0B",X"91",X"3C",
		X"80",X"0B",X"90",X"33",X"81",X"0B",X"91",X"3C",
		X"80",X"0B",X"90",X"30",X"81",X"0B",X"91",X"3C",
		X"0B",X"91",X"3F",X"0B",X"91",X"43",X"0B",X"91",
		X"3F",X"80",X"0B",X"90",X"3C",X"81",X"0B",X"90",
		X"3F",X"0B",X"90",X"3C",X"0B",X"90",X"37",X"0B",
		X"91",X"3C",X"80",X"0B",X"90",X"33",X"81",X"0B",
		X"91",X"3C",X"80",X"0B",X"90",X"30",X"81",X"0B",
		X"91",X"3C",X"0B",X"D0",X"A1",X"5C",X"5C",X"A1",
		X"5A",X"91",X"41",X"0B",X"91",X"44",X"0B",X"91",
		X"41",X"80",X"0B",X"90",X"3C",X"81",X"0B",X"90",
		X"41",X"0B",X"90",X"3C",X"0B",X"90",X"38",X"0B",
		X"91",X"3C",X"80",X"0B",X"90",X"35",X"81",X"0B",
		X"91",X"3C",X"80",X"0B",X"90",X"30",X"81",X"0B",
		X"91",X"3C",X"0B",X"91",X"41",X"0B",X"91",X"44",
		X"0B",X"91",X"41",X"80",X"0B",X"90",X"3C",X"81",
		X"0B",X"90",X"41",X"0B",X"90",X"3C",X"0B",X"90",
		X"38",X"0B",X"91",X"3C",X"80",X"0B",X"90",X"35",
		X"81",X"0B",X"91",X"3C",X"80",X"0B",X"90",X"30",
		X"81",X"0B",X"91",X"3B",X"0B",X"91",X"3E",X"0B",
		X"D0",X"A1",X"5D",X"5D",X"A1",X"5A",X"91",X"41",
		X"0B",X"91",X"3E",X"80",X"0B",X"90",X"3B",X"81",
		X"0B",X"90",X"3E",X"0B",X"90",X"3B",X"0B",X"90",
		X"38",X"0B",X"91",X"3B",X"80",X"0B",X"90",X"35",
		X"81",X"0B",X"91",X"3B",X"80",X"0B",X"90",X"30",
		X"81",X"0B",X"91",X"3B",X"0B",X"91",X"3E",X"0B",
		X"91",X"41",X"0B",X"91",X"3E",X"80",X"0B",X"90",
		X"3B",X"81",X"0B",X"90",X"3E",X"0B",X"90",X"3B",
		X"0B",X"90",X"38",X"0B",X"91",X"3B",X"80",X"0B",
		X"90",X"35",X"81",X"0B",X"91",X"3B",X"80",X"0B",
		X"90",X"30",X"81",X"0B",X"91",X"37",X"0B",X"91",
		X"3C",X"0B",X"91",X"00",X"FD",X"04",X"68",X"18",
		X"3F",X"0B",X"D0",X"A1",X"5E",X"5E",X"A1",X"5A",
		X"91",X"3C",X"80",X"0B",X"90",X"37",X"81",X"0B",
		X"90",X"3C",X"0B",X"90",X"37",X"0B",X"90",X"33",
		X"0B",X"91",X"37",X"80",X"0B",X"90",X"30",X"81",
		X"0B",X"91",X"37",X"80",X"0B",X"90",X"2E",X"81",
		X"0B",X"91",X"37",X"0B",X"91",X"3C",X"0B",X"91",
		X"3F",X"0B",X"91",X"3C",X"80",X"0B",X"90",X"37",
		X"81",X"0B",X"90",X"3C",X"0B",X"90",X"37",X"0B",
		X"90",X"33",X"0B",X"91",X"37",X"80",X"0B",X"90",
		X"30",X"81",X"0B",X"91",X"37",X"80",X"0B",X"90",
		X"2C",X"81",X"0B",X"91",X"37",X"0B",X"91",X"3C",
		X"0B",X"91",X"3F",X"0B",X"91",X"3C",X"80",X"D0",
		X"A1",X"5F",X"5F",X"A1",X"5A",X"0B",X"90",X"37",
		X"81",X"0B",X"90",X"3C",X"0B",X"90",X"37",X"0B",
		X"90",X"33",X"0B",X"91",X"37",X"80",X"0B",X"90",
		X"30",X"81",X"0B",X"91",X"37",X"80",X"0B",X"90",
		X"2B",X"81",X"0B",X"91",X"37",X"0B",X"91",X"3C",
		X"0B",X"91",X"3F",X"0B",X"91",X"3C",X"80",X"0B",
		X"90",X"37",X"81",X"0B",X"90",X"3C",X"0B",X"90",
		X"37",X"0B",X"90",X"33",X"0B",X"91",X"37",X"80",
		X"0B",X"90",X"30",X"81",X"0B",X"91",X"37",X"80",
		X"0B",X"90",X"2A",X"81",X"0B",X"91",X"39",X"0B",
		X"91",X"3C",X"0B",X"91",X"3F",X"0B",X"91",X"3C",
		X"80",X"0B",X"90",X"39",X"D0",X"A1",X"60",X"60",
		X"A1",X"5B",X"81",X"0B",X"90",X"3C",X"0B",X"90",
		X"39",X"0B",X"90",X"33",X"0B",X"91",X"39",X"80",
		X"0B",X"90",X"30",X"81",X"0B",X"91",X"39",X"80",
		X"0B",X"90",X"2A",X"81",X"0B",X"91",X"39",X"0B",
		X"91",X"3C",X"0B",X"91",X"3F",X"0B",X"91",X"3C",
		X"80",X"0B",X"90",X"39",X"81",X"0B",X"90",X"3C",
		X"0B",X"90",X"39",X"0B",X"90",X"36",X"0B",X"91",
		X"39",X"80",X"0B",X"00",X"FD",X"04",X"68",X"18",
		X"90",X"32",X"81",X"0B",X"91",X"39",X"80",X"0B",
		X"90",X"2B",X"81",X"0B",X"91",X"39",X"0B",X"91",
		X"3A",X"0B",X"91",X"3E",X"0B",X"91",X"3A",X"80",
		X"0B",X"90",X"39",X"81",X"0B",X"90",X"3A",X"D0",
		X"A1",X"61",X"61",X"A1",X"5A",X"0B",X"90",X"39",
		X"0B",X"90",X"32",X"0B",X"91",X"39",X"80",X"0B",
		X"90",X"2E",X"81",X"0B",X"91",X"39",X"80",X"0B",
		X"90",X"2B",X"81",X"0B",X"91",X"37",X"0B",X"91",
		X"3A",X"0B",X"91",X"3E",X"0B",X"91",X"3A",X"80",
		X"0B",X"90",X"37",X"81",X"0B",X"90",X"3A",X"0B",
		X"90",X"37",X"0B",X"90",X"2E",X"0B",X"91",X"37",
		X"80",X"0B",X"90",X"2B",X"81",X"0B",X"91",X"37",
		X"80",X"0B",X"90",X"27",X"81",X"0B",X"91",X"3A",
		X"0B",X"91",X"3E",X"0B",X"91",X"43",X"0B",X"91",
		X"3E",X"80",X"0B",X"90",X"3A",X"81",X"0B",X"90",
		X"3E",X"0B",X"90",X"3A",X"D0",X"A1",X"62",X"62",
		X"A1",X"5A",X"0B",X"90",X"37",X"0B",X"91",X"3A",
		X"80",X"0B",X"90",X"33",X"81",X"0B",X"91",X"3A",
		X"80",X"0B",X"90",X"30",X"81",X"0B",X"91",X"39",
		X"0B",X"91",X"3F",X"0B",X"91",X"43",X"0B",X"91",
		X"3F",X"80",X"0B",X"90",X"39",X"81",X"0B",X"90",
		X"3F",X"0B",X"90",X"39",X"0B",X"90",X"30",X"0B",
		X"91",X"39",X"80",X"0B",X"90",X"2D",X"81",X"0B",
		X"91",X"39",X"80",X"0B",X"90",X"26",X"81",X"0B",
		X"91",X"39",X"0B",X"91",X"3C",X"0B",X"91",X"42",
		X"0B",X"91",X"3C",X"80",X"0B",X"90",X"39",X"81",
		X"0B",X"90",X"3C",X"0B",X"90",X"39",X"0B",X"90",
		X"32",X"D0",X"A1",X"63",X"63",X"A1",X"5A",X"0B",
		X"91",X"39",X"80",X"0B",X"90",X"2D",X"81",X"0B",
		X"91",X"39",X"80",X"0B",X"90",X"26",X"81",X"0B",
		X"91",X"39",X"0B",X"91",X"3C",X"0B",X"91",X"42",
		X"0B",X"91",X"3C",X"00",X"FD",X"04",X"68",X"18",
		X"80",X"0B",X"90",X"39",X"81",X"0B",X"90",X"3C",
		X"0B",X"90",X"39",X"0B",X"90",X"32",X"0B",X"91",
		X"39",X"80",X"0B",X"90",X"2D",X"81",X"0B",X"91",
		X"39",X"80",X"0B",X"90",X"26",X"81",X"0B",X"91",
		X"3A",X"0B",X"91",X"3E",X"0B",X"91",X"43",X"0B",
		X"91",X"3E",X"80",X"0B",X"90",X"3A",X"81",X"0B",
		X"90",X"3E",X"0B",X"90",X"3A",X"0B",X"90",X"32",
		X"0B",X"91",X"3A",X"D0",X"A1",X"64",X"64",X"A1",
		X"59",X"80",X"0B",X"90",X"2E",X"81",X"0B",X"91",
		X"3A",X"80",X"0B",X"90",X"26",X"81",X"0B",X"91",
		X"3C",X"0B",X"91",X"42",X"0B",X"91",X"45",X"0B",
		X"91",X"42",X"80",X"0B",X"90",X"3C",X"81",X"0B",
		X"90",X"42",X"0B",X"90",X"3C",X"0B",X"90",X"33",
		X"0B",X"91",X"3C",X"80",X"0B",X"90",X"30",X"81",
		X"0B",X"91",X"3C",X"80",X"0B",X"90",X"26",X"81",
		X"0B",X"91",X"3E",X"0B",X"91",X"43",X"0B",X"91",
		X"46",X"0B",X"91",X"43",X"80",X"0B",X"90",X"3E",
		X"81",X"0B",X"90",X"43",X"0B",X"90",X"3E",X"0B",
		X"90",X"37",X"0B",X"91",X"3E",X"80",X"0B",X"D0",
		X"A1",X"65",X"65",X"A1",X"5A",X"90",X"32",X"81",
		X"0B",X"91",X"3E",X"80",X"0B",X"90",X"26",X"81",
		X"0B",X"91",X"3E",X"0B",X"91",X"42",X"0B",X"91",
		X"48",X"0B",X"91",X"42",X"80",X"0B",X"90",X"3E",
		X"81",X"0B",X"90",X"42",X"0B",X"90",X"3E",X"0B",
		X"90",X"39",X"0B",X"91",X"3E",X"80",X"0B",X"90",
		X"36",X"81",X"0B",X"91",X"3E",X"80",X"0B",X"90",
		X"26",X"81",X"0B",X"91",X"3D",X"0B",X"91",X"43",
		X"0B",X"91",X"46",X"0B",X"91",X"43",X"80",X"0B",
		X"90",X"3D",X"81",X"0B",X"90",X"43",X"0B",X"90",
		X"3D",X"0B",X"90",X"37",X"0B",X"91",X"3D",X"80",
		X"0B",X"90",X"33",X"81",X"D0",X"A1",X"66",X"66",
		X"A1",X"5A",X"0B",X"00",X"FD",X"04",X"68",X"18",
		X"91",X"3D",X"80",X"0B",X"90",X"26",X"81",X"0B",
		X"91",X"3C",X"0B",X"91",X"3F",X"0B",X"91",X"45",
		X"0B",X"91",X"3F",X"80",X"0B",X"90",X"3C",X"81",
		X"0B",X"90",X"3F",X"0B",X"90",X"3C",X"0B",X"90",
		X"36",X"0B",X"91",X"3C",X"80",X"0B",X"90",X"32",
		X"81",X"0B",X"91",X"3C",X"80",X"0B",X"90",X"26",
		X"81",X"0B",X"91",X"3A",X"0B",X"91",X"40",X"0B",
		X"91",X"43",X"0B",X"91",X"40",X"80",X"0B",X"90",
		X"3A",X"81",X"0B",X"90",X"40",X"0B",X"90",X"3A",
		X"0B",X"90",X"34",X"0B",X"91",X"3A",X"80",X"0B",
		X"90",X"31",X"81",X"0B",X"91",X"3A",X"D0",X"A1",
		X"67",X"67",X"A1",X"5B",X"80",X"0B",X"90",X"26",
		X"81",X"0B",X"91",X"39",X"0B",X"91",X"3C",X"0B",
		X"91",X"43",X"0B",X"91",X"3C",X"80",X"0B",X"90",
		X"39",X"81",X"0B",X"90",X"3C",X"0B",X"90",X"39",
		X"0B",X"90",X"33",X"0B",X"91",X"39",X"80",X"0B",
		X"90",X"30",X"81",X"0B",X"91",X"39",X"80",X"0B",
		X"90",X"26",X"81",X"0B",X"91",X"39",X"0B",X"91",
		X"3C",X"0B",X"91",X"42",X"0B",X"91",X"3C",X"80",
		X"0B",X"90",X"39",X"81",X"0B",X"90",X"3C",X"0B",
		X"90",X"39",X"0B",X"90",X"32",X"0B",X"91",X"39",
		X"80",X"0B",X"90",X"2D",X"81",X"0B",X"91",X"39",
		X"80",X"0B",X"90",X"26",X"D0",X"A1",X"68",X"68",
		X"A1",X"59",X"81",X"0B",X"91",X"37",X"0B",X"91",
		X"3A",X"0B",X"91",X"40",X"0B",X"91",X"3A",X"80",
		X"0B",X"90",X"37",X"81",X"0B",X"90",X"3A",X"0B",
		X"90",X"37",X"0B",X"90",X"31",X"0B",X"91",X"37",
		X"80",X"0B",X"90",X"2E",X"81",X"0B",X"91",X"37",
		X"80",X"0B",X"90",X"26",X"81",X"0B",X"91",X"36",
		X"0B",X"91",X"39",X"0B",X"91",X"3F",X"0B",X"91",
		X"39",X"80",X"0B",X"90",X"36",X"81",X"0B",X"90",
		X"39",X"0B",X"90",X"00",X"FD",X"04",X"68",X"18",
		X"36",X"0B",X"90",X"30",X"0B",X"91",X"36",X"80",
		X"0B",X"90",X"2D",X"81",X"0B",X"91",X"36",X"80",
		X"0B",X"90",X"26",X"81",X"0B",X"D0",X"A1",X"69",
		X"69",X"A1",X"5A",X"91",X"37",X"0B",X"91",X"3A",
		X"0B",X"91",X"3E",X"0B",X"91",X"3A",X"80",X"0B",
		X"90",X"37",X"81",X"0B",X"90",X"3A",X"0B",X"90",
		X"37",X"0B",X"90",X"2E",X"0B",X"91",X"37",X"80",
		X"0B",X"90",X"2B",X"81",X"0B",X"91",X"37",X"80",
		X"0B",X"90",X"26",X"81",X"0B",X"91",X"37",X"0B",
		X"91",X"39",X"0B",X"91",X"3C",X"0B",X"91",X"39",
		X"80",X"0B",X"90",X"37",X"81",X"0B",X"90",X"39",
		X"0B",X"90",X"37",X"0B",X"90",X"33",X"0B",X"91",
		X"37",X"80",X"0B",X"90",X"30",X"81",X"0B",X"91",
		X"37",X"80",X"0B",X"90",X"26",X"81",X"0B",X"91",
		X"36",X"0B",X"D0",X"A1",X"6A",X"6A",X"A1",X"5A",
		X"91",X"39",X"0B",X"91",X"3C",X"0B",X"91",X"39",
		X"80",X"0B",X"90",X"36",X"81",X"0B",X"90",X"39",
		X"0B",X"90",X"36",X"0B",X"90",X"32",X"0B",X"91",
		X"36",X"80",X"0B",X"90",X"2D",X"81",X"0B",X"91",
		X"36",X"80",X"0B",X"90",X"2B",X"81",X"0B",X"91",
		X"36",X"0B",X"91",X"39",X"0B",X"91",X"3C",X"0B",
		X"91",X"39",X"80",X"0B",X"90",X"36",X"81",X"0B",
		X"90",X"39",X"0B",X"90",X"36",X"0B",X"90",X"33",
		X"0B",X"91",X"36",X"80",X"0B",X"90",X"30",X"81",
		X"0B",X"91",X"36",X"80",X"0B",X"90",X"2B",X"81",
		X"0B",X"91",X"37",X"0B",X"91",X"39",X"0B",X"D0",
		X"A1",X"6B",X"6B",X"A1",X"5A",X"91",X"3C",X"0B",
		X"91",X"3B",X"80",X"0B",X"90",X"37",X"81",X"0B",
		X"90",X"3B",X"0B",X"90",X"37",X"0B",X"90",X"32",
		X"0B",X"91",X"37",X"80",X"0B",X"90",X"2F",X"81",
		X"0B",X"91",X"37",X"80",X"0B",X"90",X"2B",X"81",
		X"0B",X"91",X"39",X"00",X"FD",X"04",X"68",X"18",
		X"0B",X"91",X"3C",X"0B",X"91",X"42",X"0B",X"91",
		X"3C",X"80",X"0B",X"90",X"39",X"81",X"0B",X"90",
		X"3C",X"0B",X"90",X"39",X"0B",X"90",X"33",X"0B",
		X"91",X"39",X"80",X"0B",X"90",X"30",X"81",X"0B",
		X"91",X"39",X"80",X"0B",X"90",X"2B",X"81",X"0B",
		X"91",X"3C",X"0B",X"91",X"42",X"0B",X"91",X"45",
		X"0B",X"D0",X"A1",X"6C",X"6C",X"A1",X"5A",X"91",
		X"42",X"80",X"0B",X"90",X"3C",X"81",X"0B",X"90",
		X"42",X"0B",X"90",X"3C",X"0B",X"90",X"33",X"0B",
		X"91",X"3C",X"80",X"0B",X"90",X"30",X"81",X"0B",
		X"91",X"3C",X"80",X"0B",X"90",X"2B",X"81",X"0B",
		X"91",X"3B",X"0B",X"91",X"3E",X"0B",X"91",X"43",
		X"0B",X"91",X"3E",X"80",X"0B",X"90",X"3B",X"81",
		X"0B",X"90",X"3E",X"0B",X"90",X"3B",X"0B",X"90",
		X"37",X"0B",X"91",X"3B",X"80",X"0B",X"90",X"32",
		X"81",X"0B",X"91",X"3B",X"80",X"0B",X"90",X"2B",
		X"81",X"0B",X"91",X"3B",X"0B",X"91",X"3E",X"0B",
		X"91",X"41",X"0B",X"91",X"3E",X"80",X"D0",X"A1",
		X"6D",X"6D",X"A1",X"5A",X"0B",X"90",X"3B",X"81",
		X"0B",X"90",X"3E",X"0B",X"90",X"3B",X"0B",X"90",
		X"38",X"0B",X"91",X"3B",X"80",X"0B",X"90",X"35",
		X"81",X"0B",X"91",X"3B",X"80",X"0B",X"90",X"2B",
		X"81",X"0B",X"91",X"37",X"0B",X"91",X"3C",X"0B",
		X"91",X"3F",X"0B",X"91",X"3C",X"80",X"0B",X"90",
		X"37",X"81",X"0B",X"90",X"3C",X"0B",X"90",X"37",
		X"0B",X"90",X"33",X"0B",X"91",X"37",X"80",X"0B",
		X"90",X"30",X"81",X"0B",X"91",X"37",X"80",X"0B",
		X"90",X"2B",X"81",X"0C",X"91",X"36",X"0C",X"91",
		X"3C",X"0C",X"91",X"3F",X"0C",X"91",X"3C",X"80",
		X"0C",X"90",X"36",X"D0",X"A1",X"6E",X"6E",X"A1",
		X"5B",X"81",X"0C",X"90",X"3C",X"0C",X"90",X"36",
		X"0C",X"90",X"33",X"00",X"FD",X"04",X"68",X"18",
		X"0C",X"91",X"36",X"80",X"0C",X"90",X"30",X"81",
		X"0C",X"91",X"36",X"80",X"0C",X"90",X"2B",X"81",
		X"0C",X"91",X"36",X"0C",X"91",X"3C",X"0C",X"91",
		X"3F",X"0C",X"91",X"3C",X"80",X"0C",X"90",X"36",
		X"81",X"0C",X"90",X"3C",X"0C",X"90",X"36",X"0C",
		X"90",X"33",X"0C",X"91",X"36",X"80",X"0C",X"90",
		X"30",X"81",X"0C",X"91",X"36",X"80",X"0C",X"90",
		X"2B",X"81",X"0C",X"91",X"37",X"0C",X"91",X"3B",
		X"0C",X"91",X"3E",X"0C",X"91",X"3B",X"80",X"0D",
		X"90",X"37",X"81",X"0D",X"90",X"3B",X"D0",X"A1",
		X"6F",X"6F",X"A1",X"20",X"0D",X"90",X"3E",X"0D",
		X"90",X"3F",X"0F",X"90",X"3C",X"0F",X"90",X"39",
		X"12",X"90",X"42",X"12",X"90",X"3B",X"91",X"3E",
		X"92",X"43",X"93",X"2B",X"7F",X"80",X"81",X"82",
		X"83",X"D0",X"A1",X"70",X"70",X"A1",X"5D",X"90",
		X"45",X"91",X"36",X"0D",X"90",X"49",X"81",X"0D",
		X"91",X"42",X"90",X"4E",X"0D",X"90",X"49",X"81",
		X"0D",X"91",X"41",X"90",X"44",X"0D",X"90",X"49",
		X"81",X"0D",X"91",X"36",X"90",X"45",X"0D",X"90",
		X"49",X"81",X"0D",X"91",X"38",X"90",X"42",X"0D",
		X"90",X"49",X"81",X"0D",X"91",X"3D",X"90",X"41",
		X"0D",X"90",X"49",X"81",X"0D",X"91",X"42",X"90",
		X"45",X"0D",X"90",X"49",X"81",X"0D",X"91",X"3E",
		X"90",X"4E",X"0D",X"90",X"49",X"81",X"0D",X"91",
		X"3D",X"90",X"44",X"0D",X"90",X"49",X"81",X"0D",
		X"91",X"42",X"90",X"45",X"0D",X"90",X"49",X"81",
		X"0D",X"D0",X"A1",X"71",X"71",X"A1",X"5B",X"91",
		X"38",X"90",X"42",X"0D",X"90",X"49",X"81",X"0D",
		X"91",X"3D",X"90",X"41",X"0D",X"90",X"49",X"81",
		X"0D",X"91",X"36",X"90",X"45",X"0D",X"90",X"49",
		X"81",X"0D",X"91",X"42",X"90",X"45",X"0D",X"90",
		X"42",X"81",X"0D",X"00",X"FD",X"04",X"68",X"18",
		X"91",X"3B",X"90",X"4A",X"0D",X"90",X"47",X"81",
		X"0D",X"91",X"34",X"90",X"44",X"0D",X"90",X"47",
		X"81",X"0D",X"91",X"40",X"90",X"44",X"0D",X"90",
		X"40",X"81",X"0D",X"91",X"39",X"90",X"49",X"0D",
		X"90",X"45",X"81",X"0D",X"91",X"32",X"90",X"42",
		X"0D",X"90",X"49",X"81",X"0D",X"91",X"3E",X"90",
		X"47",X"0D",X"90",X"45",X"D0",X"A1",X"72",X"72",
		X"A1",X"59",X"81",X"0D",X"91",X"3B",X"90",X"44",
		X"0D",X"90",X"42",X"81",X"0D",X"91",X"3D",X"90",
		X"41",X"0D",X"90",X"3E",X"91",X"3D",X"0D",X"90",
		X"3D",X"91",X"41",X"0D",X"90",X"3B",X"91",X"44",
		X"0D",X"90",X"39",X"91",X"49",X"0D",X"90",X"38",
		X"91",X"47",X"0D",X"90",X"36",X"91",X"45",X"0D",
		X"90",X"49",X"81",X"0D",X"91",X"42",X"90",X"4E",
		X"0D",X"90",X"49",X"81",X"0D",X"91",X"41",X"90",
		X"44",X"0D",X"90",X"49",X"81",X"0D",X"91",X"36",
		X"90",X"45",X"0D",X"90",X"49",X"81",X"0D",X"91",
		X"38",X"90",X"42",X"0D",X"90",X"49",X"81",X"0D",
		X"D0",X"A1",X"73",X"73",X"A1",X"5B",X"91",X"3D",
		X"90",X"41",X"0D",X"90",X"49",X"81",X"0D",X"91",
		X"42",X"90",X"45",X"0D",X"90",X"49",X"81",X"0D",
		X"91",X"3E",X"90",X"4E",X"0D",X"90",X"49",X"81",
		X"0D",X"91",X"3D",X"90",X"44",X"0D",X"90",X"49",
		X"81",X"0D",X"91",X"42",X"90",X"45",X"0D",X"90",
		X"49",X"81",X"0D",X"91",X"38",X"90",X"42",X"0D",
		X"90",X"49",X"81",X"0D",X"91",X"3D",X"90",X"41",
		X"0D",X"90",X"49",X"81",X"0D",X"91",X"36",X"90",
		X"45",X"0D",X"90",X"49",X"81",X"0D",X"91",X"42",
		X"90",X"45",X"0D",X"90",X"42",X"81",X"0D",X"91",
		X"3B",X"90",X"4A",X"0D",X"90",X"47",X"D0",X"A1",
		X"74",X"74",X"A1",X"5A",X"81",X"0D",X"91",X"34",
		X"90",X"44",X"0D",X"00",X"FD",X"04",X"68",X"18",
		X"90",X"47",X"81",X"0D",X"91",X"40",X"90",X"44",
		X"0D",X"90",X"40",X"81",X"0D",X"91",X"38",X"90",
		X"4C",X"0D",X"90",X"47",X"81",X"0D",X"91",X"39",
		X"90",X"49",X"0D",X"90",X"4C",X"81",X"0D",X"91",
		X"3D",X"90",X"49",X"0D",X"90",X"45",X"81",X"0D",
		X"91",X"3D",X"90",X"40",X"0D",X"90",X"44",X"81",
		X"0D",X"91",X"39",X"90",X"45",X"0D",X"81",X"0D",
		X"91",X"34",X"0D",X"81",X"0D",X"91",X"2D",X"0D",
		X"81",X"0D",X"90",X"3D",X"91",X"4C",X"0D",X"90",
		X"40",X"91",X"4A",X"0D",X"90",X"45",X"91",X"49",
		X"D0",X"A1",X"75",X"75",X"A1",X"59",X"0D",X"90",
		X"40",X"91",X"47",X"0D",X"90",X"3B",X"91",X"45",
		X"0D",X"90",X"40",X"91",X"44",X"0D",X"90",X"3D",
		X"91",X"45",X"0D",X"90",X"40",X"91",X"47",X"0D",
		X"90",X"39",X"91",X"49",X"0D",X"90",X"40",X"91",
		X"45",X"0D",X"90",X"38",X"91",X"47",X"0D",X"90",
		X"40",X"91",X"4A",X"0D",X"90",X"39",X"91",X"49",
		X"0D",X"90",X"40",X"91",X"4A",X"0D",X"90",X"45",
		X"91",X"4C",X"0D",X"90",X"40",X"81",X"0D",X"91",
		X"44",X"90",X"3B",X"0D",X"90",X"40",X"81",X"0D",
		X"91",X"45",X"90",X"3D",X"0D",X"90",X"47",X"91",
		X"40",X"0D",X"90",X"49",X"D0",X"A1",X"76",X"76",
		X"A1",X"5A",X"91",X"39",X"0D",X"90",X"40",X"81",
		X"0D",X"91",X"47",X"90",X"38",X"0D",X"90",X"40",
		X"81",X"0D",X"91",X"49",X"90",X"3D",X"0D",X"90",
		X"40",X"81",X"0D",X"91",X"4E",X"90",X"3D",X"0D",
		X"90",X"39",X"81",X"0D",X"91",X"4B",X"90",X"42",
		X"0D",X"90",X"3F",X"81",X"0D",X"91",X"4E",X"90",
		X"3C",X"0D",X"90",X"50",X"91",X"3F",X"0D",X"90",
		X"51",X"91",X"38",X"0D",X"90",X"3F",X"81",X"0D",
		X"91",X"50",X"90",X"3C",X"0D",X"90",X"3F",X"81",
		X"0D",X"91",X"4E",X"00",X"FD",X"04",X"68",X"18",
		X"90",X"3D",X"0D",X"90",X"4C",X"81",X"0D",X"91",
		X"44",X"90",X"4B",X"0D",X"90",X"49",X"D0",X"A1",
		X"77",X"77",X"A1",X"5A",X"81",X"0D",X"91",X"38",
		X"90",X"4B",X"0D",X"90",X"48",X"81",X"0D",X"91",
		X"3D",X"90",X"49",X"0D",X"91",X"40",X"0D",X"91",
		X"44",X"0D",X"91",X"40",X"0D",X"91",X"3B",X"0D",
		X"91",X"40",X"0D",X"90",X"4C",X"91",X"3A",X"0D",
		X"91",X"3D",X"0D",X"91",X"36",X"0D",X"90",X"4E",
		X"91",X"3D",X"06",X"90",X"4F",X"06",X"90",X"3A",
		X"91",X"4E",X"0D",X"90",X"3D",X"0D",X"90",X"4C",
		X"91",X"3B",X"0D",X"90",X"4A",X"81",X"0D",X"90",
		X"4C",X"0D",X"90",X"49",X"0D",X"90",X"4A",X"0D",
		X"90",X"47",X"0D",X"91",X"3C",X"90",X"4E",X"0D",
		X"91",X"3F",X"0D",X"D0",X"A1",X"78",X"78",X"A1",
		X"5A",X"91",X"38",X"0D",X"90",X"50",X"91",X"3F",
		X"06",X"90",X"51",X"06",X"90",X"3C",X"91",X"50",
		X"0D",X"90",X"3F",X"0D",X"90",X"4E",X"91",X"3D",
		X"0D",X"90",X"4D",X"81",X"0D",X"90",X"4E",X"0D",
		X"90",X"4B",X"0D",X"90",X"4D",X"0D",X"90",X"49",
		X"0D",X"91",X"3D",X"90",X"50",X"0D",X"90",X"4D",
		X"81",X"0D",X"91",X"38",X"90",X"49",X"0D",X"90",
		X"4D",X"81",X"0D",X"91",X"35",X"90",X"50",X"0D",
		X"90",X"53",X"81",X"0D",X"91",X"31",X"90",X"56",
		X"0D",X"90",X"4D",X"81",X"0D",X"91",X"33",X"90",
		X"55",X"0D",X"90",X"4D",X"81",X"0D",X"91",X"35",
		X"D0",X"A1",X"79",X"79",X"A1",X"31",X"90",X"53",
		X"0D",X"90",X"4D",X"81",X"0D",X"91",X"39",X"90",
		X"51",X"0D",X"80",X"81",X"0D",X"90",X"3B",X"91",
		X"53",X"0D",X"90",X"51",X"81",X"0D",X"91",X"3D",
		X"90",X"50",X"0D",X"90",X"51",X"81",X"0D",X"91",
		X"36",X"90",X"4E",X"03",X"90",X"50",X"03",X"90",
		X"4E",X"47",X"80",X"00",X"FD",X"04",X"68",X"18",
		X"81",X"D0",X"A1",X"35",X"7A",X"A1",X"30",X"FF",
		X"FF",X"FF",X"15",X"15",X"FF",X"15",X"15",X"FF",
		X"FF",X"FF",X"15",X"FF",X"FF",X"FF",X"15",X"FF",
		X"15",X"FF",X"15",X"FF",X"FF",X"FF",X"15",X"FF",
		X"FF",X"FF",X"15",X"FF",X"FF",X"FF",X"15",X"FF",
		X"FF",X"FF",X"15",X"FF",X"FF",X"FF",X"15",X"FF",
		X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"7B",
		X"A1",X"30",X"FF",X"15",X"FF",X"15",X"15",X"FF",
		X"15",X"15",X"15",X"15",X"FF",X"15",X"15",X"15",
		X"FF",X"15",X"FF",X"15",X"FF",X"15",X"FF",X"15",
		X"15",X"15",X"FF",X"15",X"15",X"15",X"15",X"15",
		X"FF",X"15",X"FF",X"15",X"FF",X"15",X"FF",X"15",
		X"FF",X"15",X"FF",X"15",X"15",X"15",X"FF",X"15",
		X"FF",X"15",X"7C",X"A1",X"30",X"FF",X"15",X"FF",
		X"15",X"15",X"FF",X"15",X"15",X"FF",X"FF",X"FF",
		X"15",X"15",X"FF",X"FF",X"15",X"FF",X"FF",X"FF",
		X"15",X"FF",X"FF",X"FF",X"15",X"FF",X"FF",X"FF",
		X"15",X"15",X"15",X"FF",X"15",X"FF",X"FF",X"FF",
		X"15",X"FF",X"FF",X"FF",X"15",X"FF",X"15",X"15",
		X"15",X"15",X"FF",X"15",X"15",X"7D",X"A1",X"30",
		X"FF",X"15",X"FF",X"15",X"15",X"FF",X"15",X"15",
		X"FF",X"15",X"15",X"15",X"15",X"15",X"FF",X"15",
		X"15",X"15",X"FF",X"15",X"15",X"15",X"FF",X"15",
		X"FF",X"15",X"FF",X"15",X"15",X"15",X"FF",X"15",
		X"FF",X"15",X"FF",X"15",X"15",X"15",X"FF",X"15",
		X"FF",X"15",X"15",X"15",X"15",X"FF",X"15",X"15",
		X"7E",X"A1",X"30",X"FF",X"FF",X"FF",X"15",X"15",
		X"FF",X"15",X"15",X"FF",X"FF",X"FF",X"15",X"FF",
		X"FF",X"FF",X"15",X"15",X"15",X"FF",X"15",X"FF",
		X"FF",X"FF",X"15",X"FF",X"FF",X"FF",X"15",X"15",
		X"15",X"FF",X"15",X"FF",X"FF",X"FF",X"15",X"FF",
		X"FF",X"FF",X"15",X"00",X"FD",X"04",X"68",X"18",
		X"FF",X"FF",X"FF",X"15",X"FF",X"15",X"FF",X"15",
		X"7F",X"A1",X"07",X"06",X"30",X"30",X"30",X"30",
		X"30",X"30",X"7F",X"A8",X"07",X"06",X"30",X"30",
		X"30",X"30",X"30",X"30",X"7F",X"AF",X"03",X"02",
		X"3A",X"30",X"7F",X"B2",X"03",X"02",X"3B",X"31",
		X"00",X"00",X"54",X"65",X"74",X"72",X"6F",X"6E",
		X"69",X"73",X"F3",X"18",X"5D",X"FB",X"EE",X"19",
		X"00",X"58",X"50",X"C0",X"21",X"16",X"06",X"98",
		X"06",X"8C",X"05",X"75",X"04",X"4F",X"06",X"01",
		X"03",X"C0",X"23",X"81",X"06",X"CB",X"05",X"C0",
		X"22",X"01",X"04",X"76",X"03",X"01",X"05",X"01",
		X"06",X"B1",X"04",X"39",X"03",X"31",X"06",X"C0",
		X"20",X"1A",X"05",X"01",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"02",X"00",X"7F",X"00",X"23",X"80",
		X"FE",X"00",X"01",X"80",X"01",X"00",X"02",X"3F",
		X"3F",X"00",X"00",X"30",X"30",X"20",X"20",X"3F",
		X"2A",X"2A",X"2A",X"FC",X"01",X"FC",X"02",X"FC",
		X"03",X"FC",X"04",X"02",X"00",X"F6",X"CF",X"7E",
		X"CF",X"7C",X"11",X"00",X"50",X"2B",X"B6",X"59",
		X"00",X"2B",X"B8",X"2B",X"C6",X"CF",X"7A",X"CF",
		X"78",X"CF",X"76",X"59",X"01",X"CF",X"74",X"1A",
		X"11",X"8C",X"FF",X"82",X"03",X"35",X"3F",X"62",
		X"21",X"B8",X"35",X"72",X"27",X"59",X"F0",X"E3",
		X"10",X"2B",X"B8",X"B8",X"86",X"35",X"56",X"34",
		X"21",X"86",X"2B",X"B8",X"1A",X"11",X"82",X"01",
		X"35",X"72",X"4A",X"21",X"B6",X"99",X"B8",X"2B",
		X"B6",X"B8",X"88",X"35",X"56",X"4A",X"21",X"88",
		X"2B",X"B6",X"1A",X"11",X"82",X"02",X"35",X"72",
		X"66",X"21",X"B6",X"B8",X"B8",X"2B",X"B6",X"B8",
		X"8A",X"35",X"53",X"66",X"21",X"8A",X"2B",X"B6",
		X"90",X"66",X"59",X"00",X"2B",X"B8",X"CF",X"72",
		X"CF",X"70",X"21",X"00",X"FD",X"04",X"68",X"18",
		X"BA",X"99",X"BE",X"2B",X"C2",X"1A",X"C3",X"5E",
		X"D8",X"1A",X"BD",X"5E",X"D9",X"21",X"D8",X"AD",
		X"35",X"3F",X"8F",X"82",X"30",X"35",X"72",X"85",
		X"CF",X"6E",X"59",X"00",X"B8",X"BE",X"2B",X"BE",
		X"21",X"BA",X"2B",X"C2",X"21",X"BC",X"99",X"C0",
		X"2B",X"C4",X"1A",X"C3",X"5E",X"D8",X"1A",X"C5",
		X"5E",X"D9",X"21",X"D8",X"AD",X"35",X"3F",X"C1",
		X"82",X"30",X"35",X"72",X"AA",X"CF",X"6E",X"1A",
		X"C5",X"E6",X"6C",X"35",X"50",X"B7",X"59",X"1E",
		X"CF",X"6C",X"CF",X"6A",X"59",X"00",X"B8",X"C0",
		X"2B",X"C0",X"21",X"BC",X"2B",X"C4",X"21",X"C2",
		X"2B",X"BA",X"21",X"C4",X"2B",X"BC",X"CF",X"72",
		X"1A",X"BD",X"E6",X"7A",X"35",X"50",X"13",X"21",
		X"C8",X"35",X"3F",X"E3",X"E6",X"01",X"2B",X"C8",
		X"E3",X"23",X"CF",X"6C",X"CF",X"74",X"90",X"D2",
		X"CF",X"68",X"35",X"56",X"F0",X"CF",X"76",X"59",
		X"2A",X"CF",X"74",X"90",X"13",X"CF",X"66",X"90",
		X"02",X"03",X"00",X"E9",X"FF",X"21",X"D2",X"F3",
		X"D0",X"93",X"D0",X"93",X"D0",X"F3",X"D0",X"93",
		X"D0",X"93",X"D0",X"F3",X"D0",X"93",X"D0",X"93",
		X"D0",X"82",X"15",X"F0",X"D0",X"11",X"FA",X"00",
		X"99",X"D0",X"2B",X"D0",X"21",X"D2",X"F3",X"D0",
		X"93",X"D0",X"93",X"D0",X"F3",X"D0",X"93",X"D0",
		X"93",X"D0",X"F3",X"D0",X"93",X"D0",X"93",X"D0",
		X"82",X"2A",X"F0",X"D0",X"FF",X"75",X"59",X"07",
		X"2B",X"D6",X"59",X"0D",X"2B",X"D4",X"11",X"CE",
		X"11",X"99",X"D6",X"99",X"D6",X"F6",X"2B",X"D0",
		X"11",X"C0",X"11",X"99",X"D4",X"AD",X"99",X"D0",
		X"2B",X"D0",X"11",X"DE",X"11",X"99",X"D6",X"AD",
		X"5E",X"D2",X"5E",X"D3",X"CF",X"64",X"1A",X"D4",
		X"E6",X"01",X"5E",X"D4",X"35",X"53",X"40",X"1A",
		X"D6",X"E6",X"01",X"00",X"FD",X"04",X"68",X"18",
		X"5E",X"D6",X"35",X"53",X"3C",X"63",X"FF",X"59",
		X"76",X"5E",X"B3",X"E3",X"01",X"5E",X"B5",X"1A",
		X"B7",X"E6",X"08",X"5E",X"B2",X"5E",X"B4",X"21",
		X"96",X"F3",X"B2",X"F3",X"B4",X"93",X"B2",X"93",
		X"B2",X"93",X"B4",X"93",X"B4",X"21",X"9A",X"F3",
		X"B2",X"F3",X"B4",X"93",X"B2",X"93",X"B2",X"93",
		X"B4",X"93",X"B4",X"21",X"98",X"F3",X"B2",X"F3",
		X"B4",X"93",X"B2",X"93",X"B2",X"93",X"B4",X"93",
		X"B4",X"F3",X"B2",X"F3",X"B4",X"93",X"B2",X"93",
		X"B2",X"93",X"B4",X"93",X"B4",X"F3",X"B2",X"F3",
		X"B4",X"93",X"B2",X"93",X"B2",X"93",X"B4",X"93",
		X"B4",X"F3",X"B2",X"F3",X"B4",X"93",X"B2",X"93",
		X"B2",X"93",X"B4",X"93",X"B4",X"21",X"9A",X"F3",
		X"B2",X"F3",X"B4",X"93",X"B2",X"93",X"B2",X"93",
		X"B4",X"93",X"B4",X"21",X"96",X"F3",X"B2",X"F3",
		X"B4",X"FF",X"04",X"00",X"E0",X"FF",X"75",X"1A",
		X"D8",X"2B",X"B0",X"59",X"0D",X"2B",X"D2",X"11",
		X"C0",X"11",X"99",X"D2",X"AD",X"B8",X"B0",X"35",
		X"4D",X"68",X"E3",X"07",X"35",X"56",X"68",X"59",
		X"07",X"2B",X"D4",X"11",X"CE",X"11",X"99",X"D4",
		X"99",X"D4",X"F6",X"2B",X"D0",X"B8",X"D8",X"35",
		X"4D",X"5D",X"E3",X"FF",X"E3",X"FF",X"E3",X"02",
		X"35",X"56",X"5D",X"11",X"C0",X"11",X"99",X"D2",
		X"AD",X"99",X"D0",X"2B",X"D0",X"21",X"96",X"2B",
		X"D2",X"CF",X"64",X"CF",X"62",X"93",X"C6",X"93",
		X"C8",X"21",X"C8",X"E6",X"21",X"35",X"50",X"55",
		X"59",X"21",X"2B",X"C8",X"59",X"23",X"99",X"C8",
		X"CF",X"6C",X"63",X"FF",X"1A",X"D4",X"E6",X"01",
		X"5E",X"D4",X"35",X"53",X"1C",X"63",X"FF",X"1A",
		X"D2",X"E6",X"01",X"5E",X"D2",X"35",X"53",X"08",
		X"63",X"FF",X"59",X"14",X"5E",X"B2",X"59",X"76",
		X"5E",X"B3",X"21",X"00",X"FD",X"04",X"68",X"18",
		X"96",X"F3",X"B2",X"93",X"B3",X"F3",X"B2",X"93",
		X"B3",X"F3",X"B2",X"93",X"B3",X"F3",X"B2",X"93",
		X"B3",X"F3",X"B2",X"93",X"B3",X"F3",X"B2",X"93",
		X"B3",X"F3",X"B2",X"93",X"B3",X"F3",X"B2",X"93",
		X"B3",X"F3",X"B2",X"93",X"B3",X"F3",X"B2",X"1A",
		X"B2",X"E3",X"02",X"5E",X"B2",X"E6",X"AC",X"35",
		X"72",X"77",X"FF",X"75",X"CF",X"60",X"CF",X"70",
		X"11",X"7F",X"50",X"2B",X"BA",X"11",X"7F",X"3A",
		X"2B",X"BC",X"59",X"9A",X"2B",X"C0",X"11",X"A7",
		X"04",X"2B",X"22",X"B4",X"FD",X"35",X"4D",X"D0",
		X"FA",X"82",X"90",X"D2",X"F8",X"84",X"2B",X"BE",
		X"CF",X"5E",X"CF",X"72",X"59",X"05",X"2B",X"C8",
		X"63",X"FF",X"05",X"00",X"F6",X"FF",X"1A",X"BB",
		X"5E",X"B0",X"1A",X"BD",X"5E",X"B1",X"21",X"B0",
		X"F6",X"FC",X"9C",X"F3",X"B0",X"93",X"B1",X"21",
		X"B0",X"F6",X"FC",X"9E",X"F3",X"B0",X"FF",X"59",
		X"07",X"5E",X"B3",X"93",X"B3",X"1A",X"B3",X"5E",
		X"B5",X"E6",X"80",X"35",X"3F",X"89",X"59",X"50",
		X"5E",X"B2",X"1A",X"B3",X"E6",X"08",X"82",X"FE",
		X"35",X"3F",X"43",X"1A",X"B3",X"E6",X"18",X"82",
		X"FE",X"35",X"3F",X"43",X"21",X"96",X"2B",X"B0",
		X"90",X"49",X"21",X"94",X"2B",X"B0",X"90",X"49",
		X"59",X"A0",X"B8",X"B2",X"5E",X"B4",X"21",X"B0",
		X"F3",X"B2",X"F3",X"B4",X"93",X"B2",X"93",X"B2",
		X"1A",X"B2",X"E6",X"82",X"35",X"72",X"49",X"59",
		X"A0",X"B8",X"B2",X"5E",X"B4",X"21",X"94",X"F3",
		X"B2",X"F3",X"B4",X"93",X"B2",X"93",X"B2",X"59",
		X"A0",X"B8",X"B2",X"5E",X"B4",X"21",X"96",X"F3",
		X"B2",X"F3",X"B4",X"93",X"B2",X"93",X"B2",X"1A",
		X"B2",X"E6",X"A2",X"35",X"72",X"70",X"90",X"1C",
		X"FF",X"21",X"BE",X"35",X"53",X"A7",X"B8",X"8C",
		X"35",X"4D",X"9A",X"00",X"FD",X"04",X"68",X"18",
		X"21",X"8C",X"2B",X"BE",X"90",X"BD",X"B8",X"8E",
		X"35",X"56",X"BD",X"21",X"8C",X"99",X"8E",X"2B",
		X"BE",X"90",X"BD",X"B8",X"90",X"35",X"50",X"B2",
		X"21",X"90",X"2B",X"BE",X"90",X"BD",X"99",X"8E",
		X"35",X"53",X"BD",X"21",X"90",X"B8",X"8E",X"2B",
		X"BE",X"21",X"C0",X"B8",X"92",X"35",X"56",X"C8",
		X"21",X"92",X"2B",X"C0",X"FF",X"11",X"00",X"73",
		X"2B",X"BC",X"21",X"C2",X"B8",X"B6",X"2B",X"B0",
		X"35",X"50",X"DB",X"1A",X"B1",X"90",X"DF",X"1A",
		X"B1",X"FA",X"82",X"E9",X"2B",X"B0",X"11",X"CE",
		X"12",X"99",X"B0",X"F6",X"99",X"BE",X"2B",X"BE",
		X"21",X"C0",X"E3",X"0A",X"2B",X"C0",X"90",X"8A",
		X"06",X"00",X"F8",X"FF",X"5E",X"B0",X"1A",X"0E",
		X"B8",X"CE",X"35",X"3F",X"01",X"1A",X"0E",X"2B",
		X"CE",X"1A",X"B0",X"E6",X"01",X"35",X"72",X"FF",
		X"FF",X"75",X"11",X"C0",X"10",X"2B",X"D0",X"11",
		X"22",X"0B",X"2B",X"D2",X"CF",X"5C",X"11",X"CB",
		X"10",X"2B",X"D0",X"11",X"64",X"10",X"2B",X"D2",
		X"CF",X"5C",X"63",X"FF",X"11",X"C1",X"10",X"2B",
		X"B0",X"59",X"33",X"F0",X"B0",X"11",X"CC",X"10",
		X"2B",X"B0",X"59",X"30",X"F0",X"B0",X"93",X"B0",
		X"F0",X"B0",X"93",X"B0",X"F0",X"B0",X"93",X"B0",
		X"90",X"14",X"11",X"CE",X"10",X"2B",X"B0",X"AD",
		X"E3",X"01",X"F0",X"B0",X"E6",X"39",X"35",X"56",
		X"14",X"59",X"30",X"F0",X"B0",X"11",X"CD",X"10",
		X"2B",X"B0",X"AD",X"E3",X"01",X"F0",X"B0",X"E6",
		X"39",X"35",X"56",X"14",X"59",X"30",X"F0",X"B0",
		X"11",X"CC",X"10",X"2B",X"B0",X"AD",X"E3",X"01",
		X"F0",X"B0",X"90",X"14",X"75",X"11",X"C1",X"10",
		X"2B",X"B0",X"AD",X"E6",X"01",X"F0",X"B0",X"CF",
		X"5A",X"11",X"C1",X"10",X"2B",X"B0",X"AD",X"E6",
		X"30",X"63",X"FF",X"00",X"FD",X"04",X"68",X"18",
		X"11",X"E1",X"04",X"2B",X"22",X"59",X"00",X"5E",
		X"24",X"59",X"3F",X"5E",X"25",X"21",X"D0",X"AD",
		X"5E",X"D4",X"93",X"D0",X"21",X"D0",X"AD",X"E6",
		X"20",X"2B",X"D6",X"E9",X"E9",X"99",X"D6",X"2B",
		X"B0",X"11",X"00",X"07",X"99",X"B0",X"2B",X"B0",
		X"21",X"D6",X"E6",X"32",X"35",X"50",X"CB",X"21",
		X"B0",X"E3",X"06",X"2B",X"B0",X"59",X"05",X"5E",
		X"D5",X"21",X"D2",X"2B",X"28",X"21",X"B0",X"7F",
		X"00",X"5E",X"26",X"B4",X"CB",X"93",X"B0",X"93",
		X"D2",X"1A",X"D5",X"E6",X"01",X"5E",X"D5",X"35",
		X"72",X"CF",X"93",X"D0",X"93",X"D2",X"1A",X"D4",
		X"E6",X"01",X"5E",X"D4",X"35",X"72",X"AA",X"FF",
		X"10",X"C0",X"25",X"0A",X"33",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"03",X"30",
		X"30",X"30",X"0A",X"47",X"61",X"6D",X"65",X"20",
		X"4F",X"76",X"65",X"72",X"21",X"0A",X"59",X"6F",
		X"75",X"20",X"57",X"69",X"6E",X"21",X"21",X"21",
		X"11",X"C0",X"26",X"20",X"27",X"2E",X"35",X"3C",
		X"43",X"4A",X"51",X"58",X"5F",X"66",X"6D",X"74",
		X"7B",X"00",X"20",X"00",X"23",X"00",X"26",X"00",
		X"29",X"00",X"2C",X"00",X"2F",X"00",X"32",X"00",
		X"35",X"03",X"03",X"0B",X"0B",X"0C",X"0C",X"0F",
		X"0F",X"12",X"C0",X"1A",X"80",X"FF",X"B0",X"FF",
		X"B0",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"50",X"00",X"80",X"00",X"20",X"C0",
		X"29",X"75",X"11",X"FE",X"01",X"2B",X"B0",X"59",
		X"00",X"F3",X"B0",X"11",X"FE",X"02",X"2B",X"B0",
		X"59",X"00",X"F3",X"B0",X"11",X"FE",X"03",X"2B",
		X"B0",X"59",X"00",X"F3",X"B0",X"11",X"FE",X"04",
		X"2B",X"B0",X"59",X"00",X"F3",X"B0",X"CF",X"58",
		X"63",X"FF",X"21",X"00",X"FD",X"04",X"68",X"18",
		X"C0",X"29",X"11",X"FA",X"01",X"2B",X"B0",X"11",
		X"00",X"01",X"F3",X"B0",X"11",X"FA",X"02",X"2B",
		X"B0",X"11",X"00",X"02",X"F3",X"B0",X"11",X"FA",
		X"03",X"2B",X"B0",X"11",X"00",X"00",X"F3",X"B0",
		X"11",X"FA",X"04",X"2B",X"B0",X"11",X"00",X"00",
		X"F3",X"B0",X"FF",X"22",X"C0",X"25",X"E9",X"2B",
		X"B0",X"11",X"00",X"09",X"99",X"B0",X"2B",X"B0",
		X"7F",X"00",X"5E",X"D2",X"21",X"B0",X"7F",X"01",
		X"5E",X"D3",X"21",X"D2",X"F3",X"A0",X"F3",X"A2",
		X"59",X"00",X"F3",X"A4",X"F3",X"A6",X"59",X"03",
		X"5E",X"2C",X"FF",X"23",X"C0",X"26",X"75",X"1A",
		X"C6",X"E6",X"70",X"35",X"53",X"CB",X"11",X"CF",
		X"10",X"90",X"CE",X"11",X"DA",X"10",X"2B",X"D0",
		X"11",X"22",X"0B",X"2B",X"D2",X"CF",X"5C",X"59",
		X"01",X"CF",X"74",X"1A",X"11",X"82",X"80",X"35",
		X"72",X"D7",X"63",X"FF",X"00",X"00",X"42",X"72",
		X"69",X"63",X"6B",X"73",X"00",X"00",X"38",X"18",
		X"85",X"FB",X"EE",X"19",X"02",X"00",X"F8",X"11",
		X"DF",X"01",X"F6",X"2B",X"30",X"CD",X"C3",X"75",
		X"CF",X"32",X"35",X"50",X"10",X"CF",X"34",X"63",
		X"FF",X"21",X"36",X"AD",X"8C",X"24",X"35",X"72",
		X"21",X"11",X"CE",X"05",X"CF",X"18",X"CF",X"34",
		X"63",X"FF",X"CF",X"38",X"28",X"00",X"35",X"3F",
		X"2C",X"CF",X"3A",X"90",X"B8",X"CF",X"38",X"70",
		X"65",X"65",X"6B",X"28",X"00",X"35",X"3F",X"3E",
		X"CF",X"3A",X"AD",X"2B",X"3C",X"90",X"B8",X"CF",
		X"38",X"72",X"6E",X"64",X"28",X"00",X"35",X"3F",
		X"5C",X"CF",X"3A",X"11",X"A7",X"04",X"2B",X"22",
		X"B4",X"FD",X"35",X"50",X"4F",X"CF",X"3E",X"21",
		X"40",X"2B",X"3C",X"90",X"B8",X"CF",X"38",X"75",
		X"73",X"72",X"28",X"00",X"35",X"3F",X"6E",X"CF",
		X"3A",X"CF",X"3C",X"00",X"FD",X"04",X"68",X"18",
		X"2B",X"3C",X"90",X"B8",X"CF",X"42",X"2B",X"44",
		X"CF",X"34",X"CF",X"38",X"28",X"00",X"35",X"3F",
		X"B1",X"75",X"21",X"44",X"EC",X"00",X"CF",X"3A",
		X"35",X"53",X"87",X"CF",X"46",X"EE",X"00",X"2B",
		X"44",X"63",X"1A",X"45",X"B8",X"3C",X"E6",X"02",
		X"5E",X"45",X"21",X"48",X"FC",X"44",X"35",X"53",
		X"9F",X"21",X"48",X"90",X"A3",X"21",X"44",X"B8",
		X"48",X"35",X"53",X"A8",X"CF",X"46",X"CF",X"38",
		X"29",X"00",X"35",X"72",X"B1",X"CF",X"4A",X"21",
		X"44",X"F6",X"2B",X"3C",X"63",X"FF",X"CF",X"38",
		X"29",X"00",X"35",X"72",X"C1",X"CF",X"4A",X"63",
		X"FF",X"2B",X"4C",X"CD",X"D9",X"21",X"1A",X"2B",
		X"4E",X"21",X"4E",X"AD",X"93",X"4E",X"35",X"3F",
		X"D7",X"CF",X"50",X"90",X"CB",X"CF",X"4E",X"2B",
		X"52",X"CD",X"F1",X"1A",X"0F",X"8C",X"03",X"35",
		X"72",X"F0",X"21",X"54",X"2B",X"50",X"CF",X"56",
		X"42",X"72",X"65",X"61",X"6B",X"00",X"FF",X"2B",
		X"58",X"93",X"1B",X"FF",X"03",X"00",X"F9",X"CD",
		X"6E",X"2B",X"44",X"E6",X"83",X"35",X"4D",X"6D",
		X"1A",X"31",X"E6",X"78",X"35",X"4D",X"6D",X"1A",
		X"30",X"E6",X"9A",X"35",X"56",X"19",X"75",X"CF",
		X"5A",X"63",X"21",X"44",X"E6",X"52",X"35",X"53",
		X"29",X"E3",X"32",X"2B",X"40",X"11",X"00",X"07",
		X"90",X"2E",X"2B",X"40",X"11",X"00",X"08",X"2B",
		X"44",X"21",X"40",X"35",X"50",X"6D",X"E9",X"E9",
		X"99",X"40",X"99",X"44",X"2B",X"44",X"11",X"E1",
		X"04",X"2B",X"22",X"21",X"2A",X"2B",X"24",X"21",
		X"30",X"2B",X"28",X"EC",X"FE",X"E3",X"06",X"2B",
		X"30",X"59",X"05",X"2B",X"40",X"21",X"44",X"7F",
		X"00",X"5E",X"26",X"B4",X"CB",X"93",X"44",X"93",
		X"28",X"21",X"40",X"E6",X"01",X"35",X"4D",X"52",
		X"5E",X"26",X"B4",X"00",X"FD",X"04",X"68",X"18",
		X"CB",X"EE",X"FE",X"FF",X"2B",X"50",X"2B",X"54",
		X"CD",X"F4",X"75",X"2B",X"4E",X"11",X"00",X"0B",
		X"2B",X"22",X"1A",X"21",X"E6",X"38",X"35",X"50",
		X"87",X"E6",X"FF",X"B4",X"E6",X"11",X"A0",X"1B",
		X"2B",X"36",X"21",X"4E",X"F3",X"36",X"59",X"A2",
		X"5E",X"36",X"59",X"7F",X"CF",X"50",X"2B",X"30",
		X"1A",X"0F",X"2B",X"4E",X"1A",X"0F",X"F0",X"36",
		X"FC",X"4E",X"35",X"72",X"AC",X"21",X"36",X"AD",
		X"90",X"9C",X"21",X"36",X"AD",X"8C",X"0A",X"35",
		X"3F",X"EF",X"8C",X"75",X"35",X"72",X"D0",X"59",
		X"20",X"CF",X"50",X"2B",X"30",X"1A",X"30",X"E6",
		X"06",X"35",X"50",X"CE",X"5E",X"30",X"21",X"36",
		X"E6",X"01",X"2B",X"36",X"90",X"94",X"E6",X"60",
		X"35",X"53",X"94",X"1A",X"30",X"E6",X"96",X"35",
		X"50",X"E6",X"59",X"A2",X"5E",X"36",X"59",X"5C",
		X"CF",X"50",X"90",X"94",X"21",X"36",X"AD",X"CF",
		X"50",X"93",X"36",X"90",X"94",X"11",X"E8",X"06",
		X"CF",X"18",X"93",X"1B",X"FF",X"04",X"00",X"F8",
		X"2B",X"5C",X"CD",X"EF",X"CF",X"34",X"CF",X"38",
		X"67",X"6F",X"74",X"6F",X"00",X"35",X"3F",X"12",
		X"CF",X"3A",X"CF",X"5E",X"CF",X"38",X"67",X"6F",
		X"73",X"75",X"62",X"00",X"35",X"3F",X"26",X"CF",
		X"3A",X"75",X"21",X"36",X"EC",X"00",X"CF",X"5E",
		X"CF",X"38",X"72",X"65",X"74",X"75",X"72",X"6E",
		X"00",X"35",X"3F",X"3F",X"1A",X"1C",X"35",X"72",
		X"39",X"CF",X"60",X"F6",X"2B",X"36",X"63",X"CF",
		X"62",X"CF",X"38",X"69",X"66",X"00",X"35",X"3F",
		X"96",X"CF",X"3A",X"DF",X"FC",X"EC",X"02",X"CF",
		X"64",X"35",X"72",X"54",X"CF",X"4A",X"EC",X"00",
		X"CF",X"3A",X"CF",X"38",X"74",X"68",X"65",X"6E",
		X"00",X"EE",X"02",X"FC",X"3C",X"35",X"53",X"6A",
		X"EE",X"02",X"90",X"00",X"FD",X"04",X"68",X"18",
		X"6E",X"EE",X"02",X"B8",X"3C",X"35",X"56",X"73",
		X"59",X"04",X"35",X"53",X"78",X"59",X"01",X"35",
		X"72",X"7D",X"59",X"02",X"2B",X"40",X"EE",X"00",
		X"F8",X"40",X"DF",X"04",X"35",X"3F",X"8A",X"CF",
		X"66",X"21",X"36",X"AD",X"35",X"3F",X"94",X"93",
		X"36",X"90",X"8A",X"CF",X"62",X"CF",X"38",X"70",
		X"6F",X"6B",X"65",X"00",X"35",X"3F",X"B3",X"CF",
		X"3A",X"2B",X"68",X"CF",X"38",X"2C",X"00",X"35",
		X"72",X"AD",X"CF",X"4A",X"CF",X"3A",X"F0",X"68",
		X"CF",X"62",X"CF",X"38",X"27",X"00",X"35",X"72",
		X"C0",X"CF",X"38",X"72",X"65",X"6D",X"00",X"35",
		X"3F",X"CF",X"21",X"36",X"AD",X"35",X"3F",X"CD",
		X"93",X"36",X"90",X"C3",X"CF",X"62",X"CF",X"38",
		X"6C",X"69",X"6E",X"65",X"00",X"35",X"3F",X"DE",
		X"11",X"A0",X"19",X"CF",X"18",X"CF",X"38",X"65",
		X"6E",X"64",X"00",X"35",X"3F",X"EA",X"CF",X"56",
		X"00",X"11",X"00",X"05",X"CF",X"18",X"2B",X"66",
		X"93",X"1B",X"93",X"1B",X"FF",X"05",X"00",X"00",
		X"CF",X"38",X"6E",X"65",X"78",X"74",X"00",X"35",
		X"3F",X"37",X"CF",X"42",X"2B",X"68",X"75",X"21",
		X"36",X"EC",X"00",X"11",X"00",X"FF",X"99",X"68",
		X"F6",X"35",X"72",X"1C",X"CF",X"46",X"2B",X"36",
		X"CF",X"3A",X"21",X"68",X"F6",X"E3",X"01",X"F3",
		X"68",X"B8",X"3C",X"35",X"56",X"32",X"EE",X"00",
		X"2B",X"36",X"CF",X"34",X"63",X"CF",X"58",X"CF",
		X"62",X"CF",X"38",X"66",X"6F",X"72",X"00",X"35",
		X"3F",X"6C",X"CF",X"42",X"2B",X"68",X"CF",X"34",
		X"CF",X"38",X"3D",X"00",X"35",X"72",X"4F",X"CF",
		X"4A",X"CF",X"3A",X"F3",X"68",X"CF",X"38",X"74",
		X"6F",X"00",X"35",X"72",X"5D",X"CF",X"4A",X"11",
		X"00",X"FF",X"99",X"68",X"2B",X"6A",X"21",X"36",
		X"F3",X"6A",X"CF",X"00",X"FD",X"04",X"68",X"18",
		X"3A",X"CF",X"62",X"CF",X"38",X"61",X"74",X"00",
		X"35",X"3F",X"9A",X"CF",X"3A",X"35",X"53",X"7B",
		X"CF",X"46",X"5E",X"30",X"CF",X"38",X"2C",X"00",
		X"35",X"3F",X"98",X"CF",X"3A",X"35",X"53",X"8B",
		X"CF",X"46",X"E6",X"78",X"35",X"50",X"92",X"CF",
		X"46",X"E3",X"F8",X"E9",X"AD",X"5E",X"31",X"CF",
		X"62",X"CF",X"38",X"70",X"75",X"74",X"00",X"35",
		X"3F",X"A9",X"CF",X"3A",X"CF",X"50",X"CF",X"62",
		X"CF",X"38",X"6D",X"6F",X"64",X"65",X"00",X"35",
		X"3F",X"C7",X"CF",X"3A",X"1A",X"21",X"E6",X"20",
		X"35",X"50",X"C5",X"11",X"00",X"0B",X"2B",X"22",
		X"21",X"3C",X"B4",X"E6",X"CF",X"62",X"11",X"A0",
		X"14",X"CF",X"18",X"59",X"00",X"2B",X"3C",X"E9",
		X"E9",X"E9",X"E9",X"2B",X"40",X"93",X"36",X"21",
		X"36",X"AD",X"E6",X"30",X"35",X"50",X"FD",X"E6",
		X"0A",X"35",X"53",X"EB",X"E3",X"0A",X"99",X"40",
		X"90",X"CE",X"82",X"DF",X"E6",X"07",X"35",X"50",
		X"FD",X"E6",X"06",X"35",X"53",X"FD",X"E3",X"10",
		X"99",X"40",X"90",X"CE",X"FF",X"06",X"00",X"FD",
		X"CD",X"BB",X"75",X"CF",X"32",X"35",X"56",X"B9",
		X"21",X"48",X"2B",X"40",X"2B",X"6A",X"FC",X"6C",
		X"35",X"3F",X"16",X"21",X"48",X"CF",X"6E",X"F6",
		X"B8",X"3C",X"35",X"50",X"5A",X"21",X"6C",X"2B",
		X"40",X"21",X"40",X"F6",X"B8",X"3C",X"35",X"53",
		X"2D",X"21",X"40",X"CF",X"70",X"90",X"1D",X"35",
		X"56",X"5A",X"21",X"00",X"FC",X"48",X"35",X"3F",
		X"58",X"21",X"6A",X"2B",X"44",X"CF",X"6E",X"2B",
		X"6A",X"2B",X"4E",X"21",X"4E",X"AD",X"F0",X"44",
		X"93",X"4E",X"93",X"44",X"21",X"4E",X"82",X"1F",
		X"35",X"72",X"41",X"21",X"6A",X"FC",X"40",X"35",
		X"72",X"37",X"59",X"01",X"35",X"3F",X"70",X"21",
		X"00",X"E6",X"80",X"00",X"FD",X"04",X"68",X"18",
		X"E6",X"C0",X"FC",X"48",X"35",X"72",X"6A",X"CF",
		X"4A",X"21",X"48",X"CF",X"70",X"2B",X"48",X"21",
		X"36",X"AD",X"35",X"3F",X"8A",X"21",X"3C",X"F3",
		X"40",X"93",X"40",X"93",X"40",X"21",X"36",X"AD",
		X"93",X"36",X"F0",X"40",X"35",X"72",X"7C",X"90",
		X"B7",X"21",X"40",X"2B",X"6A",X"FC",X"48",X"35",
		X"3F",X"B1",X"21",X"6A",X"CF",X"70",X"2B",X"6A",
		X"2B",X"4E",X"21",X"4E",X"AD",X"F0",X"40",X"93",
		X"4E",X"93",X"40",X"21",X"4E",X"82",X"1F",X"35",
		X"72",X"9B",X"21",X"6A",X"2B",X"40",X"90",X"8E",
		X"21",X"48",X"CF",X"6E",X"2B",X"48",X"21",X"3C",
		X"63",X"FF",X"2B",X"72",X"11",X"3F",X"35",X"2B",
		X"2A",X"11",X"A0",X"18",X"2B",X"5A",X"CF",X"18",
		X"CF",X"52",X"2A",X"2A",X"2A",X"20",X"54",X"69",
		X"6E",X"79",X"20",X"42",X"41",X"53",X"49",X"43",
		X"20",X"44",X"45",X"56",X"00",X"CF",X"5A",X"11",
		X"A0",X"08",X"2B",X"1A",X"FF",X"59",X"00",X"F0",
		X"36",X"59",X"20",X"CF",X"50",X"CF",X"5A",X"59",
		X"A2",X"5E",X"36",X"CF",X"34",X"21",X"36",X"AD",
		X"63",X"FF",X"08",X"A0",X"5F",X"CD",X"B6",X"88",
		X"1F",X"E3",X"01",X"2B",X"4E",X"35",X"56",X"B3",
		X"82",X"E0",X"35",X"72",X"B3",X"21",X"4E",X"E3",
		X"A0",X"FF",X"21",X"4E",X"FF",X"2B",X"70",X"CD",
		X"CE",X"E6",X"20",X"2B",X"4E",X"35",X"50",X"CB",
		X"82",X"60",X"35",X"72",X"CB",X"21",X"4E",X"E6",
		X"A0",X"FF",X"21",X"4E",X"FF",X"2B",X"6E",X"CD",
		X"FA",X"21",X"6C",X"2B",X"40",X"FC",X"48",X"35",
		X"3F",X"F3",X"21",X"40",X"F6",X"FC",X"3C",X"35",
		X"72",X"ED",X"21",X"40",X"E3",X"02",X"2B",X"36",
		X"CF",X"58",X"CF",X"66",X"21",X"40",X"CF",X"70",
		X"90",X"D4",X"CF",X"56",X"4C",X"69",X"6E",X"65",
		X"00",X"93",X"1B",X"00",X"FD",X"04",X"68",X"18",
		X"FF",X"09",X"A0",X"5E",X"2B",X"5E",X"CD",X"DE",
		X"75",X"35",X"53",X"B0",X"59",X"00",X"B8",X"3C",
		X"2B",X"3C",X"59",X"2D",X"CF",X"50",X"59",X"00",
		X"2B",X"44",X"21",X"3C",X"35",X"53",X"C4",X"11",
		X"D0",X"8A",X"99",X"3C",X"2B",X"3C",X"59",X"03",
		X"2B",X"44",X"11",X"10",X"27",X"CF",X"74",X"11",
		X"E8",X"03",X"CF",X"74",X"59",X"64",X"CF",X"74",
		X"59",X"0A",X"CF",X"74",X"59",X"30",X"99",X"3C",
		X"CF",X"50",X"63",X"FF",X"2B",X"76",X"CD",X"EA",
		X"CF",X"56",X"53",X"74",X"61",X"63",X"6B",X"00",
		X"2B",X"60",X"CD",X"F7",X"CF",X"56",X"53",X"79",
		X"6E",X"74",X"61",X"78",X"00",X"2B",X"4A",X"93",
		X"1B",X"FF",X"0A",X"A0",X"5F",X"CD",X"D2",X"21",
		X"1A",X"2B",X"4E",X"21",X"36",X"2B",X"6A",X"21",
		X"4E",X"AD",X"93",X"4E",X"35",X"3F",X"CE",X"2B",
		X"40",X"21",X"36",X"AD",X"88",X"20",X"FC",X"40",
		X"35",X"72",X"C0",X"93",X"36",X"90",X"A8",X"21",
		X"6A",X"2B",X"36",X"21",X"4E",X"AD",X"93",X"4E",
		X"35",X"72",X"C4",X"CF",X"4E",X"CF",X"34",X"CF",
		X"4E",X"2B",X"38",X"CD",X"FA",X"11",X"00",X"80",
		X"2B",X"3C",X"E9",X"E9",X"99",X"3C",X"E9",X"2B",
		X"40",X"21",X"36",X"AD",X"E6",X"30",X"35",X"50",
		X"F7",X"E6",X"0A",X"35",X"53",X"F7",X"E3",X"0A",
		X"99",X"40",X"93",X"36",X"90",X"D9",X"21",X"3C",
		X"FF",X"93",X"1B",X"FF",X"0B",X"A0",X"60",X"2B",
		X"32",X"CD",X"D1",X"21",X"36",X"AD",X"35",X"3F",
		X"B3",X"8C",X"3A",X"35",X"72",X"B1",X"93",X"36",
		X"CF",X"66",X"CF",X"4A",X"21",X"36",X"CF",X"70",
		X"2B",X"36",X"FC",X"48",X"35",X"3F",X"CE",X"11",
		X"C0",X"1B",X"FC",X"36",X"35",X"3F",X"CE",X"21",
		X"36",X"E3",X"02",X"2B",X"36",X"CF",X"66",X"CF",
		X"56",X"00",X"2B",X"00",X"FD",X"04",X"68",X"18",
		X"62",X"CD",X"FB",X"21",X"00",X"2B",X"40",X"59",
		X"02",X"2B",X"6A",X"21",X"40",X"E6",X"36",X"2B",
		X"40",X"59",X"00",X"F0",X"40",X"93",X"40",X"1A",
		X"40",X"35",X"72",X"E3",X"21",X"6A",X"E6",X"01",
		X"35",X"72",X"DB",X"11",X"C0",X"1B",X"2B",X"6C",
		X"FF",X"93",X"1B",X"FF",X"0C",X"A0",X"60",X"2B",
		X"78",X"CD",X"ED",X"75",X"1A",X"1C",X"E6",X"8D",
		X"35",X"53",X"AC",X"CF",X"60",X"CF",X"38",X"2D",
		X"00",X"35",X"3F",X"BB",X"CF",X"7A",X"59",X"00",
		X"B8",X"3C",X"90",X"C1",X"CF",X"38",X"2B",X"00",
		X"CF",X"7A",X"75",X"EC",X"00",X"CF",X"38",X"2B",
		X"00",X"35",X"3F",X"D5",X"CF",X"7A",X"EE",X"00",
		X"99",X"3C",X"EC",X"00",X"90",X"C4",X"CF",X"38",
		X"2D",X"00",X"35",X"3F",X"E6",X"CF",X"7A",X"EE",
		X"00",X"B8",X"3C",X"EC",X"00",X"90",X"C4",X"EE",
		X"00",X"2B",X"3C",X"63",X"63",X"FF",X"2B",X"3A",
		X"CD",X"F9",X"CF",X"56",X"56",X"61",X"6C",X"75",
		X"65",X"00",X"2B",X"46",X"93",X"1B",X"FF",X"0D",
		X"A0",X"60",X"CD",X"E4",X"75",X"CF",X"4C",X"75",
		X"21",X"3C",X"EC",X"00",X"CF",X"38",X"2A",X"00",
		X"35",X"3F",X"B9",X"CF",X"4C",X"EE",X"00",X"CF",
		X"7C",X"EC",X"00",X"90",X"A8",X"CF",X"38",X"2F",
		X"00",X"35",X"3F",X"CA",X"CF",X"4C",X"EE",X"00",
		X"CF",X"3E",X"EC",X"00",X"90",X"A8",X"CF",X"38",
		X"25",X"00",X"35",X"3F",X"DD",X"CF",X"4C",X"EE",
		X"00",X"CF",X"3E",X"21",X"40",X"EC",X"00",X"90",
		X"A8",X"EE",X"00",X"2B",X"3C",X"63",X"63",X"FF",
		X"2B",X"7A",X"93",X"1B",X"FF",X"CF",X"38",X"72",
		X"75",X"6E",X"00",X"35",X"3F",X"F9",X"CF",X"78",
		X"F6",X"2B",X"3C",X"CF",X"5E",X"11",X"A0",X"16",
		X"CF",X"18",X"0E",X"A0",X"60",X"CD",X"FB",X"2B",
		X"6A",X"FC",X"3C",X"00",X"FD",X"04",X"68",X"18",
		X"2B",X"44",X"21",X"6A",X"35",X"53",X"B1",X"59",
		X"00",X"B8",X"6A",X"2B",X"6A",X"21",X"3C",X"35",
		X"53",X"BC",X"59",X"00",X"B8",X"3C",X"2B",X"3C",
		X"35",X"72",X"C1",X"CF",X"46",X"59",X"00",X"2B",
		X"40",X"2B",X"4E",X"21",X"40",X"99",X"40",X"2B",
		X"40",X"21",X"6A",X"35",X"53",X"D4",X"93",X"40",
		X"21",X"6A",X"99",X"6A",X"2B",X"6A",X"21",X"40",
		X"B8",X"3C",X"35",X"50",X"E5",X"2B",X"40",X"93",
		X"6A",X"21",X"4E",X"E3",X"01",X"82",X"0F",X"35",
		X"72",X"C5",X"21",X"44",X"35",X"53",X"F8",X"59",
		X"00",X"B8",X"6A",X"FF",X"21",X"6A",X"FF",X"93",
		X"1B",X"FF",X"0F",X"A0",X"5E",X"2B",X"3E",X"CD",
		X"C7",X"2B",X"4E",X"59",X"00",X"2B",X"6A",X"59",
		X"01",X"2B",X"40",X"F8",X"4E",X"35",X"3F",X"B7",
		X"21",X"6A",X"99",X"3C",X"2B",X"6A",X"21",X"3C",
		X"99",X"3C",X"2B",X"3C",X"21",X"40",X"99",X"40",
		X"35",X"72",X"AA",X"21",X"6A",X"FF",X"2B",X"7C",
		X"CD",X"E6",X"21",X"00",X"2B",X"40",X"21",X"36",
		X"AD",X"82",X"5F",X"E6",X"40",X"35",X"50",X"E4",
		X"E6",X"1B",X"35",X"53",X"E4",X"93",X"36",X"E9",
		X"99",X"40",X"FF",X"CF",X"4A",X"2B",X"42",X"CD",
		X"F7",X"21",X"36",X"AD",X"8C",X"20",X"35",X"72",
		X"F6",X"93",X"36",X"90",X"EA",X"FF",X"2B",X"34",
		X"93",X"1B",X"FF",X"10",X"A0",X"60",X"CD",X"FB",
		X"75",X"21",X"6C",X"2B",X"6A",X"FC",X"48",X"35",
		X"3F",X"C9",X"CF",X"58",X"21",X"6A",X"F6",X"2B",
		X"3C",X"CF",X"76",X"93",X"6A",X"93",X"6A",X"21",
		X"6A",X"AD",X"35",X"3F",X"C1",X"CF",X"50",X"90",
		X"B5",X"CF",X"5A",X"21",X"6A",X"CF",X"70",X"90",
		X"A3",X"2B",X"3C",X"21",X"00",X"E6",X"80",X"E6",
		X"C0",X"FC",X"6A",X"35",X"3F",X"E2",X"21",X"6A",
		X"CF",X"70",X"2B",X"00",X"FD",X"04",X"68",X"18",
		X"6A",X"21",X"3C",X"E3",X"20",X"90",X"C9",X"21",
		X"50",X"FC",X"54",X"35",X"72",X"F9",X"CF",X"76",
		X"CF",X"52",X"20",X"62",X"79",X"74",X"65",X"73",
		X"20",X"66",X"72",X"65",X"65",X"00",X"63",X"FF",
		X"93",X"1B",X"FF",X"11",X"A0",X"60",X"2B",X"7E",
		X"CD",X"C1",X"75",X"2B",X"40",X"21",X"3C",X"B8",
		X"40",X"35",X"50",X"B2",X"2B",X"3C",X"93",X"44",
		X"90",X"A7",X"21",X"44",X"35",X"3F",X"BF",X"88",
		X"30",X"CF",X"50",X"59",X"30",X"2B",X"44",X"63",
		X"FF",X"2B",X"74",X"CD",X"F1",X"75",X"59",X"00",
		X"2B",X"44",X"CF",X"38",X"3C",X"00",X"35",X"3F",
		X"D3",X"93",X"44",X"CF",X"38",X"3E",X"00",X"35",
		X"3F",X"E0",X"21",X"44",X"E3",X"04",X"2B",X"44",
		X"CF",X"38",X"3D",X"00",X"35",X"3F",X"ED",X"21",
		X"44",X"E3",X"02",X"2B",X"44",X"21",X"44",X"63",
		X"FF",X"2B",X"64",X"11",X"A0",X"1B",X"F6",X"2B",
		X"48",X"E3",X"02",X"93",X"1B",X"FF",X"12",X"A0",
		X"5D",X"2B",X"36",X"CD",X"F7",X"21",X"1A",X"2B",
		X"4E",X"1A",X"30",X"E6",X"02",X"35",X"56",X"AF",
		X"CF",X"5A",X"59",X"00",X"5E",X"1C",X"21",X"4E",
		X"AD",X"35",X"3F",X"E3",X"59",X"3F",X"CF",X"50",
		X"21",X"4E",X"AD",X"93",X"4E",X"35",X"72",X"BB",
		X"CF",X"52",X"20",X"65",X"72",X"72",X"6F",X"72",
		X"00",X"E6",X"20",X"F8",X"36",X"F6",X"35",X"3F",
		X"E1",X"2B",X"3C",X"CF",X"52",X"20",X"69",X"6E",
		X"20",X"00",X"CF",X"76",X"CF",X"5A",X"CF",X"52",
		X"4F",X"6B",X"00",X"CF",X"5A",X"59",X"00",X"CF",
		X"5C",X"35",X"3F",X"EA",X"CF",X"72",X"35",X"4D",
		X"EA",X"11",X"2B",X"56",X"CF",X"66",X"13",X"A0",
		X"59",X"21",X"36",X"AD",X"35",X"3F",X"F3",X"8C",
		X"3A",X"35",X"3F",X"F3",X"21",X"36",X"AD",X"35",
		X"3F",X"F1",X"8C",X"00",X"FD",X"04",X"68",X"18",
		X"3A",X"35",X"3F",X"F1",X"8C",X"18",X"35",X"72",
		X"CE",X"93",X"36",X"CF",X"38",X"22",X"00",X"35",
		X"72",X"CC",X"21",X"36",X"AD",X"35",X"3F",X"CC",
		X"CF",X"50",X"90",X"B9",X"90",X"D2",X"CF",X"3A",
		X"CF",X"76",X"CF",X"38",X"2C",X"00",X"35",X"3F",
		X"E8",X"59",X"20",X"CF",X"50",X"1A",X"30",X"E6",
		X"02",X"82",X"07",X"35",X"72",X"D9",X"90",X"A9",
		X"CF",X"38",X"3B",X"00",X"35",X"72",X"A9",X"CF",
		X"5A",X"90",X"F5",X"CF",X"5A",X"CF",X"62",X"14",
		X"A0",X"5F",X"CF",X"38",X"3F",X"00",X"35",X"72",
		X"AD",X"CF",X"38",X"70",X"72",X"69",X"6E",X"74",
		X"00",X"35",X"3F",X"B5",X"11",X"A0",X"13",X"CF",
		X"18",X"CF",X"38",X"69",X"6E",X"70",X"75",X"74",
		X"00",X"35",X"3F",X"F8",X"21",X"36",X"AD",X"CF",
		X"50",X"CF",X"42",X"2B",X"68",X"CF",X"34",X"DF",
		X"FC",X"21",X"36",X"EC",X"02",X"88",X"1F",X"E6",
		X"1F",X"F6",X"EC",X"00",X"59",X"3F",X"CF",X"50",
		X"CF",X"5A",X"EE",X"00",X"CF",X"5C",X"35",X"3F",
		X"D8",X"CF",X"3A",X"F3",X"68",X"EE",X"02",X"2B",
		X"36",X"DF",X"04",X"CF",X"38",X"2C",X"00",X"35",
		X"72",X"C0",X"CF",X"62",X"11",X"A0",X"15",X"CF",
		X"18",X"15",X"A0",X"58",X"CF",X"38",X"63",X"6C",
		X"73",X"00",X"35",X"3F",X"CB",X"11",X"00",X"01",
		X"AD",X"5E",X"31",X"59",X"0E",X"2B",X"6A",X"CF",
		X"5A",X"21",X"6A",X"E6",X"01",X"35",X"4D",X"AF",
		X"CF",X"5A",X"11",X"00",X"01",X"AD",X"8C",X"08",
		X"35",X"72",X"BA",X"59",X"08",X"5E",X"31",X"CF",
		X"62",X"CF",X"38",X"6C",X"69",X"73",X"74",X"00",
		X"35",X"3F",X"D9",X"CF",X"7E",X"CF",X"62",X"CF",
		X"38",X"73",X"61",X"76",X"65",X"00",X"35",X"3F",
		X"F1",X"1A",X"21",X"E6",X"28",X"35",X"53",X"EC",
		X"CF",X"46",X"11",X"00",X"FD",X"04",X"68",X"18",
		X"A0",X"17",X"CF",X"18",X"11",X"EB",X"0D",X"CF",
		X"18",X"16",X"A0",X"60",X"CF",X"38",X"6E",X"65",
		X"77",X"00",X"35",X"3F",X"B0",X"CF",X"78",X"2B",
		X"48",X"CF",X"7E",X"CF",X"56",X"00",X"CF",X"38",
		X"6C",X"65",X"74",X"00",X"CF",X"42",X"2B",X"68",
		X"CF",X"34",X"CF",X"38",X"28",X"00",X"35",X"3F",
		X"EF",X"CF",X"3A",X"35",X"53",X"CA",X"CF",X"46",
		X"1A",X"69",X"B8",X"3C",X"E6",X"02",X"5E",X"69",
		X"21",X"48",X"FC",X"68",X"35",X"53",X"DD",X"21",
		X"48",X"90",X"E1",X"21",X"68",X"B8",X"48",X"35",
		X"53",X"E6",X"CF",X"46",X"CF",X"38",X"29",X"00",
		X"35",X"72",X"EF",X"CF",X"4A",X"CF",X"38",X"3D",
		X"00",X"35",X"72",X"F8",X"CF",X"4A",X"CF",X"3A",
		X"F3",X"68",X"CF",X"62",X"17",X"A0",X"5F",X"21",
		X"00",X"5E",X"27",X"E6",X"60",X"2B",X"68",X"CD",
		X"E8",X"75",X"2B",X"44",X"1A",X"27",X"E3",X"08",
		X"5E",X"27",X"1A",X"30",X"E6",X"06",X"35",X"53",
		X"DE",X"59",X"0A",X"F0",X"68",X"21",X"68",X"88",
		X"1F",X"8C",X"1F",X"2B",X"68",X"2B",X"24",X"59",
		X"01",X"5E",X"26",X"11",X"06",X"0B",X"2B",X"22",
		X"B4",X"E6",X"35",X"3F",X"DA",X"59",X"03",X"5E",
		X"0F",X"CF",X"58",X"59",X"08",X"5E",X"27",X"21",
		X"44",X"F0",X"68",X"93",X"68",X"CF",X"54",X"63",
		X"FF",X"2B",X"50",X"1A",X"0F",X"8C",X"FF",X"35",
		X"72",X"EA",X"CF",X"7E",X"59",X"20",X"CF",X"50",
		X"21",X"54",X"2B",X"50",X"CF",X"62",X"18",X"A0",
		X"60",X"11",X"E1",X"04",X"2B",X"22",X"59",X"00",
		X"5E",X"30",X"5E",X"26",X"1A",X"31",X"E3",X"0F",
		X"82",X"78",X"35",X"72",X"B4",X"59",X"08",X"5E",
		X"31",X"21",X"2A",X"2B",X"24",X"21",X"30",X"2B",
		X"28",X"B4",X"CB",X"93",X"28",X"B4",X"CB",X"93",
		X"28",X"1A",X"28",X"00",X"FD",X"04",X"68",X"18",
		X"8C",X"A0",X"35",X"72",X"BE",X"11",X"00",X"01",
		X"2B",X"40",X"88",X"FF",X"F6",X"B8",X"30",X"1A",
		X"19",X"35",X"72",X"F9",X"21",X"40",X"E3",X"10",
		X"2B",X"24",X"AD",X"5E",X"26",X"21",X"40",X"AD",
		X"F0",X"24",X"1A",X"26",X"F0",X"40",X"93",X"40",
		X"93",X"40",X"1A",X"40",X"8C",X"E0",X"35",X"72",
		X"DC",X"93",X"30",X"93",X"30",X"FF",X"19",X"A0",
		X"60",X"59",X"01",X"2B",X"24",X"11",X"00",X"01",
		X"2B",X"26",X"CF",X"3A",X"75",X"EC",X"00",X"CF",
		X"38",X"2C",X"00",X"35",X"72",X"B5",X"CF",X"4A",
		X"CF",X"3A",X"2B",X"6A",X"35",X"53",X"C8",X"59",
		X"00",X"B8",X"26",X"2B",X"26",X"59",X"00",X"B8",
		X"6A",X"2B",X"6A",X"EE",X"00",X"2B",X"40",X"35",
		X"53",X"DB",X"59",X"00",X"B8",X"24",X"2B",X"24",
		X"59",X"00",X"B8",X"40",X"2B",X"40",X"B8",X"6A",
		X"35",X"53",X"F8",X"21",X"40",X"2B",X"4E",X"21",
		X"6A",X"2B",X"40",X"21",X"4E",X"2B",X"6A",X"21",
		X"24",X"2B",X"4E",X"21",X"26",X"2B",X"24",X"21",
		X"4E",X"2B",X"26",X"63",X"11",X"A0",X"1A",X"CF",
		X"18",X"1A",X"A0",X"60",X"21",X"3C",X"35",X"53",
		X"A8",X"11",X"00",X"78",X"90",X"AB",X"11",X"00",
		X"88",X"2B",X"28",X"21",X"40",X"2B",X"4E",X"2B",
		X"44",X"1A",X"2B",X"F0",X"30",X"21",X"4E",X"E6",
		X"01",X"2B",X"4E",X"35",X"50",X"FC",X"21",X"44",
		X"B8",X"6A",X"B8",X"6A",X"2B",X"44",X"35",X"53",
		X"D7",X"99",X"40",X"99",X"40",X"2B",X"44",X"21",
		X"26",X"99",X"30",X"2B",X"30",X"21",X"24",X"99",
		X"30",X"2B",X"30",X"1A",X"30",X"E6",X"A0",X"35",
		X"50",X"ED",X"35",X"56",X"EB",X"93",X"31",X"E3",
		X"40",X"5E",X"30",X"1A",X"31",X"82",X"78",X"35",
		X"72",X"FA",X"21",X"28",X"99",X"30",X"2B",X"30",
		X"90",X"B3",X"CF",X"00",X"FD",X"04",X"68",X"18",
		X"62",X"1B",X"A0",X"06",X"A0",X"1B",X"4E",X"45",
		X"57",X"00",X"00",X"54",X"69",X"6E",X"79",X"42",
		X"41",X"53",X"49",X"8C",X"18",X"8B",X"FB",X"EE",
		X"19",X"02",X"00",X"10",X"59",X"AD",X"2B",X"22",
		X"11",X"A0",X"FF",X"2B",X"1A",X"11",X"8C",X"8B",
		X"2B",X"24",X"B4",X"E2",X"FF",X"A0",X"0C",X"11",
		X"00",X"02",X"2B",X"1A",X"11",X"3C",X"98",X"2B",
		X"24",X"B4",X"E2",X"00",X"1B",X"C0",X"19",X"64",
		X"00",X"27",X"54",X"49",X"43",X"2D",X"54",X"41",
		X"43",X"2D",X"54",X"4F",X"45",X"2E",X"20",X"59",
		X"4F",X"55",X"20",X"28",X"58",X"29",X"20",X"00",
		X"1B",X"E0",X"15",X"D2",X"00",X"3F",X"22",X"54",
		X"4F",X"4D",X"20",X"50",X"49",X"54",X"54",X"4D",
		X"41",X"4E",X"27",X"53",X"20",X"22",X"3B",X"00",
		X"1C",X"A0",X"12",X"D3",X"00",X"3F",X"22",X"54",
		X"49",X"43",X"2D",X"54",X"41",X"43",X"2D",X"54",
		X"4F",X"45",X"2E",X"22",X"00",X"1C",X"C0",X"12",
		X"D4",X"00",X"3F",X"22",X"59",X"4F",X"55",X"20",
		X"41",X"47",X"41",X"49",X"4E",X"53",X"54",X"22",
		X"3B",X"00",X"1C",X"E0",X"11",X"D5",X"00",X"3F",
		X"22",X"20",X"54",X"49",X"4E",X"59",X"20",X"42",
		X"41",X"53",X"49",X"43",X"22",X"00",X"1D",X"A0",
		X"16",X"DD",X"00",X"3F",X"22",X"59",X"4F",X"55",
		X"20",X"41",X"52",X"45",X"20",X"58",X"2E",X"20",
		X"49",X"20",X"41",X"4D",X"22",X"3B",X"00",X"1D",
		X"C0",X"0D",X"DE",X"00",X"3F",X"22",X"20",X"4F",
		X"2E",X"20",X"59",X"4F",X"55",X"22",X"00",X"1D",
		X"E0",X"10",X"E7",X"00",X"3F",X"22",X"50",X"4C",
		X"41",X"59",X"20",X"59",X"4F",X"55",X"52",X"22",
		X"3B",X"00",X"1E",X"A0",X"15",X"E8",X"00",X"3F",
		X"22",X"20",X"54",X"55",X"52",X"4E",X"20",X"42",
		X"59",X"20",X"54",X"00",X"FD",X"04",X"68",X"18",
		X"59",X"50",X"49",X"4E",X"47",X"22",X"00",X"1E",
		X"C0",X"16",X"E9",X"00",X"3F",X"22",X"54",X"48",
		X"45",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",
		X"20",X"4F",X"46",X"20",X"41",X"22",X"3B",X"00",
		X"1E",X"E0",X"0E",X"EA",X"00",X"3F",X"22",X"20",
		X"53",X"51",X"55",X"41",X"52",X"45",X"2E",X"22",
		X"00",X"1F",X"A0",X"06",X"F0",X"00",X"41",X"3D",
		X"30",X"00",X"1F",X"C0",X"06",X"FA",X"00",X"42",
		X"3D",X"30",X"00",X"1F",X"E0",X"06",X"04",X"01",
		X"43",X"3D",X"30",X"00",X"20",X"A0",X"06",X"0E",
		X"01",X"44",X"3D",X"30",X"00",X"20",X"C0",X"06",
		X"18",X"01",X"45",X"3D",X"30",X"00",X"20",X"E0",
		X"06",X"22",X"01",X"46",X"3D",X"30",X"00",X"21",
		X"A0",X"06",X"E8",X"03",X"46",X"3D",X"31",X"00",
		X"21",X"C0",X"04",X"F2",X"03",X"3F",X"00",X"21",
		X"E0",X"0F",X"FC",X"03",X"3F",X"22",X"4E",X"45",
		X"57",X"20",X"47",X"41",X"4D",X"45",X"2E",X"22",
		X"00",X"22",X"A0",X"06",X"4C",X"04",X"49",X"3D",
		X"37",X"00",X"22",X"C0",X"0F",X"56",X"04",X"41",
		X"28",X"49",X"29",X"3D",X"30",X"3A",X"49",X"3D",
		X"49",X"2B",X"31",X"00",X"22",X"E0",X"11",X"60",
		X"04",X"49",X"46",X"49",X"3C",X"31",X"36",X"47",
		X"4F",X"54",X"4F",X"31",X"31",X"31",X"30",X"00",
		X"23",X"A0",X"06",X"6A",X"04",X"55",X"3D",X"39",
		X"00",X"23",X"C0",X"06",X"74",X"04",X"5A",X"3D",
		X"30",X"00",X"23",X"E0",X"10",X"7F",X"04",X"49",
		X"46",X"46",X"3D",X"30",X"47",X"4F",X"54",X"4F",
		X"34",X"30",X"31",X"30",X"00",X"24",X"A0",X"0B",
		X"89",X"04",X"47",X"4F",X"54",X"4F",X"32",X"30",
		X"31",X"30",X"00",X"24",X"C0",X"06",X"E6",X"05",
		X"5A",X"3D",X"31",X"00",X"24",X"E0",X"06",X"F0",
		X"05",X"46",X"3D",X"00",X"FD",X"04",X"68",X"18",
		X"30",X"00",X"25",X"A0",X"06",X"DA",X"07",X"49",
		X"3D",X"36",X"00",X"25",X"C0",X"08",X"3E",X"08",
		X"49",X"3D",X"49",X"2B",X"31",X"00",X"25",X"E0",
		X"08",X"48",X"08",X"3F",X"22",X"20",X"22",X"3B",
		X"00",X"26",X"A0",X"13",X"53",X"08",X"47",X"4F",
		X"54",X"4F",X"41",X"28",X"49",X"29",X"2A",X"32",
		X"30",X"2B",X"32",X"32",X"30",X"30",X"00",X"26",
		X"C0",X"08",X"98",X"08",X"3F",X"49",X"2D",X"36",
		X"3B",X"00",X"26",X"E0",X"0B",X"A2",X"08",X"47",
		X"4F",X"54",X"4F",X"32",X"33",X"30",X"30",X"00",
		X"27",X"A0",X"08",X"AC",X"08",X"3F",X"22",X"58",
		X"22",X"3B",X"00",X"27",X"C0",X"0B",X"B6",X"08",
		X"47",X"4F",X"54",X"4F",X"32",X"33",X"30",X"30",
		X"00",X"27",X"E0",X"08",X"D4",X"08",X"3F",X"22",
		X"4F",X"22",X"3B",X"00",X"28",X"A0",X"14",X"FC",
		X"08",X"49",X"46",X"49",X"2F",X"33",X"2A",X"33",
		X"3D",X"49",X"47",X"4F",X"54",X"4F",X"32",X"34",
		X"30",X"30",X"00",X"28",X"C0",X"09",X"06",X"09",
		X"3F",X"22",X"20",X"7C",X"22",X"3B",X"00",X"28",
		X"E0",X"0B",X"10",X"09",X"47",X"4F",X"54",X"4F",
		X"32",X"31",X"31",X"30",X"00",X"29",X"A0",X"04",
		X"60",X"09",X"3F",X"00",X"29",X"C0",X"11",X"74",
		X"09",X"49",X"46",X"49",X"3D",X"31",X"35",X"47",
		X"4F",X"54",X"4F",X"33",X"30",X"30",X"30",X"00",
		X"29",X"E0",X"11",X"7E",X"09",X"3F",X"22",X"2D",
		X"2D",X"2D",X"2B",X"2D",X"2D",X"2D",X"2B",X"2D",
		X"2D",X"2D",X"22",X"00",X"2A",X"A0",X"0B",X"88",
		X"09",X"47",X"4F",X"54",X"4F",X"32",X"31",X"31",
		X"30",X"00",X"2A",X"C0",X"10",X"B8",X"0B",X"49",
		X"46",X"5A",X"3D",X"30",X"47",X"4F",X"54",X"4F",
		X"33",X"31",X"30",X"30",X"00",X"2A",X"E0",X"10",
		X"CC",X"0B",X"49",X"00",X"FD",X"04",X"68",X"18",
		X"46",X"46",X"3D",X"31",X"47",X"4F",X"54",X"4F",
		X"33",X"30",X"35",X"30",X"00",X"2B",X"A0",X"0E",
		X"D6",X"0B",X"3F",X"22",X"59",X"4F",X"55",X"20",
		X"57",X"49",X"4E",X"2E",X"22",X"00",X"2B",X"C0",
		X"0B",X"E0",X"0B",X"47",X"4F",X"54",X"4F",X"31",
		X"30",X"31",X"30",X"00",X"2B",X"E0",X"0C",X"EA",
		X"0B",X"3F",X"22",X"49",X"20",X"57",X"49",X"4E",
		X"2E",X"22",X"00",X"2C",X"A0",X"0B",X"F4",X"0B",
		X"47",X"4F",X"54",X"4F",X"31",X"30",X"31",X"30",
		X"00",X"2C",X"C0",X"10",X"1C",X"0C",X"49",X"46",
		X"55",X"3E",X"30",X"47",X"4F",X"54",X"4F",X"33",
		X"32",X"31",X"30",X"00",X"2C",X"E0",X"11",X"26",
		X"0C",X"3F",X"22",X"43",X"41",X"54",X"27",X"53",
		X"20",X"47",X"41",X"4D",X"45",X"2E",X"22",X"00",
		X"2D",X"A0",X"08",X"30",X"0C",X"46",X"3D",X"31",
		X"2D",X"46",X"00",X"2D",X"C0",X"0B",X"3A",X"0C",
		X"47",X"4F",X"54",X"4F",X"31",X"30",X"31",X"30",
		X"00",X"2D",X"E0",X"0F",X"8A",X"0C",X"3F",X"22",
		X"59",X"4F",X"55",X"52",X"20",X"50",X"4C",X"41",
		X"22",X"3B",X"00",X"2E",X"A0",X"0D",X"97",X"0C",
		X"49",X"4E",X"50",X"55",X"54",X"59",X"3A",X"49",
		X"3D",X"59",X"00",X"2E",X"C0",X"11",X"9F",X"0C",
		X"49",X"46",X"49",X"3C",X"3D",X"30",X"47",X"4F",
		X"54",X"4F",X"33",X"32",X"34",X"30",X"00",X"2E",
		X"E0",X"11",X"A0",X"0C",X"49",X"46",X"49",X"3C",
		X"31",X"30",X"47",X"4F",X"54",X"4F",X"33",X"32",
		X"37",X"30",X"00",X"2F",X"A0",X"14",X"A8",X"0C",
		X"3F",X"22",X"50",X"4C",X"45",X"41",X"53",X"45",
		X"20",X"54",X"59",X"50",X"45",X"20",X"41",X"22",
		X"3B",X"00",X"2F",X"C0",X"0D",X"AA",X"0C",X"3F",
		X"22",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",
		X"22",X"00",X"2F",X"00",X"FD",X"04",X"68",X"18",
		X"E0",X"16",X"AB",X"0C",X"3F",X"22",X"42",X"45",
		X"54",X"57",X"45",X"45",X"4E",X"20",X"31",X"20",
		X"41",X"4E",X"44",X"20",X"39",X"22",X"3B",X"00",
		X"30",X"A0",X"10",X"B3",X"0C",X"3F",X"22",X"20",
		X"57",X"48",X"45",X"52",X"45",X"20",X"59",X"4F",
		X"55",X"22",X"00",X"30",X"C0",X"13",X"B4",X"0C",
		X"3F",X"22",X"57",X"49",X"53",X"48",X"20",X"54",
		X"4F",X"20",X"50",X"4C",X"41",X"59",X"22",X"3B",
		X"00",X"30",X"E0",X"0D",X"B5",X"0C",X"3F",X"22",
		X"20",X"59",X"4F",X"55",X"52",X"20",X"58",X"22",
		X"00",X"31",X"A0",X"0B",X"BC",X"0C",X"47",X"4F",
		X"54",X"4F",X"33",X"32",X"31",X"30",X"00",X"31",
		X"C0",X"15",X"C6",X"0C",X"49",X"46",X"41",X"28",
		X"49",X"2B",X"36",X"29",X"3D",X"30",X"47",X"4F",
		X"54",X"4F",X"33",X"33",X"31",X"30",X"00",X"31",
		X"E0",X"15",X"D1",X"0C",X"3F",X"22",X"54",X"48",
		X"41",X"54",X"20",X"53",X"51",X"55",X"41",X"52",
		X"45",X"20",X"49",X"53",X"22",X"3B",X"00",X"32",
		X"A0",X"17",X"D2",X"0C",X"3F",X"22",X"20",X"41",
		X"4C",X"52",X"45",X"41",X"44",X"59",X"22",X"3A",
		X"3F",X"22",X"54",X"41",X"4B",X"45",X"4E",X"22",
		X"00",X"32",X"C0",X"0B",X"DA",X"0C",X"47",X"4F",
		X"54",X"4F",X"33",X"32",X"31",X"30",X"00",X"32",
		X"E0",X"11",X"EE",X"0C",X"41",X"28",X"49",X"2B",
		X"36",X"29",X"3D",X"31",X"3A",X"55",X"3D",X"55",
		X"2D",X"31",X"00",X"33",X"A0",X"09",X"F8",X"0C",
		X"57",X"3D",X"36",X"31",X"30",X"30",X"00",X"33",
		X"C0",X"09",X"02",X"0D",X"47",X"4F",X"53",X"55",
		X"42",X"57",X"00",X"33",X"E0",X"11",X"0D",X"0D",
		X"49",X"46",X"4A",X"3C",X"3D",X"30",X"47",X"4F",
		X"54",X"4F",X"33",X"33",X"35",X"30",X"00",X"34",
		X"A0",X"14",X"0E",X"00",X"FD",X"04",X"68",X"18",
		X"0D",X"49",X"46",X"4C",X"2A",X"4D",X"2A",X"4E",
		X"3D",X"31",X"47",X"4F",X"54",X"4F",X"31",X"35",
		X"31",X"30",X"00",X"34",X"C0",X"0A",X"16",X"0D",
		X"57",X"3D",X"57",X"2B",X"31",X"30",X"30",X"00",
		X"34",X"E0",X"13",X"20",X"0D",X"49",X"46",X"57",
		X"3C",X"36",X"35",X"30",X"30",X"47",X"4F",X"54",
		X"4F",X"33",X"33",X"33",X"30",X"00",X"35",X"A0",
		X"10",X"52",X"0D",X"49",X"46",X"55",X"3D",X"30",
		X"47",X"4F",X"54",X"4F",X"32",X"30",X"31",X"30",
		X"00",X"35",X"C0",X"06",X"AA",X"0F",X"49",X"3D",
		X"31",X"00",X"35",X"E0",X"07",X"B4",X"0F",X"54",
		X"3D",X"2D",X"31",X"00",X"36",X"A0",X"06",X"CC",
		X"10",X"53",X"3D",X"30",X"00",X"36",X"C0",X"15",
		X"D7",X"10",X"49",X"46",X"41",X"28",X"49",X"2B",
		X"36",X"29",X"3E",X"30",X"47",X"4F",X"54",X"4F",
		X"34",X"34",X"38",X"30",X"00",X"36",X"E0",X"09",
		X"E0",X"10",X"57",X"3D",X"36",X"31",X"30",X"30",
		X"00",X"37",X"A0",X"09",X"EA",X"10",X"47",X"4F",
		X"53",X"55",X"42",X"57",X"00",X"37",X"C0",X"10",
		X"F4",X"10",X"49",X"46",X"4A",X"3D",X"30",X"47",
		X"4F",X"54",X"4F",X"34",X"34",X"31",X"30",X"00",
		X"37",X"E0",X"0A",X"FE",X"10",X"4A",X"3D",X"4C",
		X"2B",X"4D",X"2B",X"4E",X"00",X"38",X"A0",X"10",
		X"09",X"11",X"49",X"46",X"4A",X"3D",X"34",X"47",
		X"4F",X"54",X"4F",X"34",X"34",X"31",X"30",X"00",
		X"38",X"C0",X"0E",X"13",X"11",X"49",X"46",X"4A",
		X"3D",X"32",X"53",X"3D",X"53",X"2B",X"32",X"30",
		X"00",X"38",X"E0",X"0F",X"1D",X"11",X"49",X"46",
		X"4A",X"3D",X"36",X"53",X"3D",X"53",X"2B",X"31",
		X"30",X"30",X"00",X"39",X"A0",X"0D",X"27",X"11",
		X"49",X"46",X"4A",X"3D",X"30",X"53",X"3D",X"53",
		X"2B",X"32",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"39",X"C0",X"08",X"30",X"11",X"53",X"3D",X"53",
		X"2B",X"4A",X"00",X"39",X"E0",X"0A",X"3A",X"11",
		X"57",X"3D",X"57",X"2B",X"31",X"30",X"30",X"00",
		X"3A",X"A0",X"13",X"44",X"11",X"49",X"46",X"57",
		X"3C",X"36",X"35",X"30",X"30",X"47",X"4F",X"54",
		X"4F",X"34",X"33",X"33",X"30",X"00",X"3A",X"C0",
		X"10",X"4F",X"11",X"49",X"46",X"53",X"3C",X"54",
		X"47",X"4F",X"54",X"4F",X"34",X"34",X"37",X"30",
		X"00",X"3A",X"E0",X"06",X"58",X"11",X"54",X"3D",
		X"53",X"00",X"3B",X"A0",X"06",X"62",X"11",X"42",
		X"3D",X"49",X"00",X"3B",X"C0",X"08",X"76",X"11",
		X"3F",X"22",X"2E",X"22",X"3B",X"00",X"3B",X"E0",
		X"08",X"80",X"11",X"49",X"3D",X"49",X"2B",X"31",
		X"00",X"3C",X"A0",X"11",X"8A",X"11",X"49",X"46",
		X"49",X"3C",X"31",X"30",X"47",X"4F",X"54",X"4F",
		X"34",X"33",X"30",X"30",X"00",X"3C",X"C0",X"0F",
		X"94",X"11",X"3F",X"22",X"49",X"20",X"50",X"4C",
		X"41",X"59",X"20",X"22",X"3B",X"42",X"00",X"3C",
		X"E0",X"04",X"9E",X"11",X"3F",X"00",X"3D",X"A0",
		X"0B",X"A9",X"11",X"41",X"28",X"42",X"2B",X"36",
		X"29",X"3D",X"33",X"00",X"3D",X"C0",X"08",X"B2",
		X"11",X"55",X"3D",X"55",X"2D",X"31",X"00",X"3D",
		X"E0",X"12",X"BD",X"11",X"49",X"46",X"54",X"3C",
		X"31",X"30",X"30",X"47",X"4F",X"54",X"4F",X"32",
		X"30",X"31",X"30",X"00",X"3E",X"A0",X"06",X"D0",
		X"11",X"46",X"3D",X"31",X"00",X"3E",X"C0",X"06",
		X"DA",X"11",X"5A",X"3D",X"31",X"00",X"3E",X"E0",
		X"0B",X"E4",X"11",X"47",X"4F",X"54",X"4F",X"32",
		X"30",X"31",X"30",X"00",X"3F",X"A0",X"10",X"D4",
		X"17",X"4A",X"3D",X"28",X"49",X"2D",X"31",X"29",
		X"2F",X"33",X"2A",X"33",X"2B",X"38",X"00",X"3F",
		X"C0",X"06",X"DE",X"00",X"FD",X"04",X"68",X"18",
		X"17",X"44",X"3D",X"31",X"00",X"3F",X"E0",X"0B",
		X"E8",X"17",X"47",X"4F",X"54",X"4F",X"36",X"35",
		X"30",X"30",X"00",X"40",X"A0",X"12",X"38",X"18",
		X"4A",X"3D",X"49",X"2D",X"28",X"49",X"2D",X"31",
		X"29",X"2F",X"33",X"2A",X"33",X"2B",X"39",X"00",
		X"40",X"C0",X"06",X"42",X"18",X"44",X"3D",X"33",
		X"00",X"40",X"E0",X"0B",X"4C",X"18",X"47",X"4F",
		X"54",X"4F",X"36",X"35",X"30",X"30",X"00",X"41",
		X"A0",X"13",X"9C",X"18",X"49",X"46",X"49",X"25",
		X"34",X"3C",X"3E",X"31",X"47",X"4F",X"54",X"4F",
		X"36",X"34",X"34",X"30",X"00",X"41",X"C0",X"06",
		X"A6",X"18",X"44",X"3D",X"34",X"00",X"41",X"E0",
		X"07",X"BA",X"18",X"4A",X"3D",X"31",X"31",X"00",
		X"42",X"A0",X"0B",X"C4",X"18",X"47",X"4F",X"54",
		X"4F",X"36",X"35",X"30",X"30",X"00",X"42",X"C0",
		X"06",X"00",X"19",X"44",X"3D",X"32",X"00",X"42",
		X"E0",X"11",X"0B",X"19",X"49",X"46",X"49",X"3C",
		X"3D",X"31",X"47",X"4F",X"54",X"4F",X"36",X"34",
		X"34",X"30",X"00",X"43",X"A0",X"11",X"0C",X"19",
		X"49",X"46",X"49",X"3E",X"3D",X"39",X"47",X"4F",
		X"54",X"4F",X"36",X"34",X"34",X"30",X"00",X"43",
		X"C0",X"12",X"0D",X"19",X"49",X"46",X"49",X"25",
		X"32",X"3D",X"31",X"47",X"4F",X"54",X"4F",X"36",
		X"33",X"33",X"30",X"00",X"43",X"E0",X"06",X"28",
		X"19",X"4A",X"3D",X"30",X"00",X"44",X"A0",X"09",
		X"32",X"19",X"52",X"45",X"54",X"55",X"52",X"4E",
		X"00",X"44",X"C0",X"0B",X"64",X"19",X"4C",X"3D",
		X"41",X"28",X"4A",X"2D",X"44",X"29",X"00",X"44",
		X"E0",X"09",X"66",X"19",X"4D",X"3D",X"41",X"28",
		X"4A",X"29",X"00",X"45",X"A0",X"0B",X"6E",X"19",
		X"4E",X"3D",X"41",X"28",X"4A",X"2B",X"44",X"29",
		X"00",X"45",X"C0",X"00",X"FD",X"04",X"68",X"18",
		X"09",X"82",X"19",X"52",X"45",X"54",X"55",X"52",
		X"4E",X"00",X"45",X"E2",X"04",X"52",X"55",X"4E",
		X"00",X"1B",X"A0",X"02",X"E0",X"45",X"00",X"00",
		X"54",X"69",X"63",X"54",X"61",X"63",X"00",X"00",
		X"19",X"18",X"98",X"FB",X"EE",X"19",X"02",X"00",
		X"E2",X"CD",X"0A",X"2A",X"2A",X"20",X"57",X"6F",
		X"7A",X"4D",X"6F",X"6E",X"00",X"2B",X"30",X"11",
		X"DF",X"01",X"F6",X"2B",X"32",X"CD",X"60",X"E6",
		X"52",X"35",X"53",X"22",X"E3",X"32",X"2B",X"34",
		X"11",X"00",X"07",X"90",X"27",X"2B",X"34",X"11",
		X"00",X"08",X"2B",X"36",X"21",X"34",X"E9",X"E9",
		X"99",X"34",X"99",X"36",X"2B",X"36",X"11",X"E1",
		X"04",X"2B",X"22",X"21",X"2A",X"2B",X"24",X"21",
		X"32",X"2B",X"28",X"EC",X"FE",X"E3",X"06",X"2B",
		X"32",X"59",X"05",X"2B",X"34",X"21",X"36",X"7F",
		X"00",X"5E",X"26",X"B4",X"CB",X"93",X"36",X"93",
		X"28",X"21",X"34",X"E6",X"01",X"35",X"4D",X"48",
		X"EE",X"FE",X"FF",X"2B",X"38",X"CD",X"AD",X"1A",
		X"32",X"35",X"3F",X"AC",X"11",X"E1",X"04",X"2B",
		X"22",X"11",X"00",X"08",X"5E",X"32",X"99",X"32",
		X"35",X"53",X"7B",X"11",X"00",X"08",X"2B",X"32",
		X"2B",X"28",X"5E",X"26",X"B4",X"CB",X"93",X"28",
		X"1A",X"28",X"8C",X"A0",X"35",X"72",X"81",X"11",
		X"EE",X"01",X"2B",X"34",X"21",X"34",X"AD",X"E6",
		X"78",X"35",X"53",X"9D",X"8C",X"80",X"90",X"9F",
		X"8C",X"08",X"F0",X"34",X"21",X"34",X"E6",X"02",
		X"2B",X"34",X"8C",X"FE",X"35",X"72",X"91",X"FF",
		X"2B",X"3A",X"CD",X"D9",X"75",X"2B",X"30",X"11",
		X"52",X"06",X"2B",X"22",X"21",X"30",X"B4",X"F5",
		X"E6",X"0A",X"35",X"50",X"C4",X"E3",X"07",X"E3",
		X"3A",X"CF",X"38",X"21",X"30",X"82",X"0F",X"E6",
		X"0A",X"35",X"50",X"00",X"FD",X"04",X"68",X"18",
		X"D3",X"E3",X"07",X"E3",X"3A",X"CF",X"38",X"63",
		X"FF",X"2B",X"3C",X"11",X"00",X"03",X"CF",X"18",
		X"03",X"00",X"F3",X"CD",X"D3",X"75",X"59",X"80",
		X"2B",X"3E",X"CF",X"3A",X"93",X"3E",X"21",X"3E",
		X"AD",X"35",X"3F",X"D1",X"E6",X"2E",X"35",X"50",
		X"07",X"35",X"72",X"1D",X"59",X"01",X"2B",X"40",
		X"90",X"07",X"E6",X"0C",X"35",X"72",X"28",X"E6",
		X"01",X"2B",X"40",X"90",X"07",X"E6",X"18",X"35",
		X"72",X"31",X"CF",X"42",X"90",X"07",X"59",X"00",
		X"2B",X"30",X"2B",X"44",X"E9",X"E9",X"E9",X"E9",
		X"2B",X"34",X"21",X"3E",X"AD",X"93",X"3E",X"E6",
		X"30",X"35",X"50",X"68",X"E6",X"0A",X"35",X"53",
		X"54",X"2B",X"30",X"E3",X"0A",X"99",X"34",X"90",
		X"35",X"E6",X"06",X"82",X"1F",X"35",X"56",X"68",
		X"E6",X"07",X"35",X"53",X"68",X"2B",X"30",X"E3",
		X"10",X"99",X"34",X"90",X"35",X"21",X"30",X"35",
		X"3F",X"CD",X"21",X"3E",X"E6",X"02",X"2B",X"3E",
		X"21",X"40",X"35",X"53",X"84",X"21",X"44",X"F0",
		X"46",X"21",X"46",X"E3",X"01",X"2B",X"46",X"90",
		X"07",X"35",X"72",X"91",X"CF",X"3A",X"21",X"44",
		X"2B",X"46",X"E6",X"01",X"2B",X"42",X"21",X"42",
		X"B8",X"44",X"35",X"53",X"C7",X"21",X"42",X"E3",
		X"01",X"2B",X"42",X"82",X"07",X"35",X"72",X"A5",
		X"CF",X"3A",X"1A",X"32",X"35",X"72",X"BA",X"59",
		X"02",X"5E",X"32",X"1A",X"43",X"CF",X"3C",X"1A",
		X"42",X"CF",X"3C",X"59",X"3A",X"CF",X"38",X"21",
		X"32",X"E3",X"04",X"2B",X"32",X"21",X"42",X"AD",
		X"CF",X"3C",X"90",X"91",X"59",X"00",X"2B",X"40",
		X"90",X"07",X"59",X"5C",X"CF",X"38",X"63",X"FF",
		X"2B",X"48",X"93",X"32",X"11",X"20",X"0F",X"2B",
		X"2A",X"5E",X"24",X"CF",X"3A",X"59",X"2A",X"CF",
		X"38",X"21",X"30",X"00",X"FD",X"04",X"68",X"18",
		X"AD",X"93",X"30",X"35",X"72",X"E2",X"11",X"00",
		X"04",X"CF",X"18",X"04",X"00",X"72",X"59",X"81",
		X"2B",X"3E",X"CF",X"3A",X"59",X"7F",X"5E",X"2B",
		X"CF",X"38",X"2B",X"32",X"1A",X"0F",X"2B",X"30",
		X"1A",X"0F",X"F0",X"3E",X"FC",X"30",X"35",X"72",
		X"1E",X"21",X"3E",X"AD",X"90",X"0E",X"21",X"3E",
		X"AD",X"8C",X"0A",X"35",X"3F",X"60",X"8C",X"75",
		X"35",X"72",X"42",X"59",X"20",X"CF",X"38",X"2B",
		X"32",X"1A",X"32",X"E6",X"06",X"35",X"50",X"40",
		X"5E",X"32",X"21",X"3E",X"E6",X"01",X"2B",X"3E",
		X"90",X"04",X"E6",X"60",X"35",X"53",X"04",X"1A",
		X"32",X"8C",X"96",X"35",X"72",X"57",X"59",X"5C",
		X"CF",X"38",X"11",X"00",X"04",X"CF",X"18",X"21",
		X"3E",X"AD",X"CF",X"38",X"93",X"3E",X"90",X"04",
		X"F0",X"3E",X"2B",X"40",X"59",X"20",X"CF",X"38",
		X"59",X"0F",X"5E",X"2B",X"CF",X"48",X"90",X"FE",
		X"00",X"57",X"6F",X"7A",X"4D",X"6F",X"6E",X"00",
		X"00",X"26",X"18",X"A0",X"FB",X"EE",X"19",X"02",
		X"00",X"54",X"1A",X"21",X"E6",X"40",X"35",X"53",
		X"0B",X"21",X"0E",X"F3",X"17",X"90",X"05",X"59",
		X"A0",X"2B",X"24",X"11",X"60",X"7E",X"2B",X"26",
		X"11",X"03",X"0B",X"2B",X"22",X"B4",X"F3",X"11",
		X"EE",X"01",X"2B",X"7A",X"59",X"7E",X"F0",X"7A",
		X"1A",X"7A",X"E6",X"02",X"5E",X"7A",X"35",X"53",
		X"20",X"11",X"01",X"01",X"2B",X"7A",X"59",X"60",
		X"F0",X"7A",X"11",X"FF",X"10",X"2B",X"7A",X"11",
		X"F6",X"01",X"2B",X"7C",X"11",X"00",X"5E",X"F3",
		X"7C",X"59",X"FE",X"5E",X"0E",X"11",X"00",X"5F",
		X"2B",X"1A",X"11",X"AC",X"5E",X"FF",X"03",X"00",
		X"CF",X"A2",X"24",X"BD",X"93",X"03",X"20",X"EF",
		X"FF",X"CA",X"D0",X"F7",X"86",X"E2",X"E6",X"E3",
		X"D0",X"02",X"E6",X"00",X"FD",X"04",X"68",X"18",
		X"E4",X"AD",X"11",X"D0",X"10",X"F5",X"20",X"C6",
		X"03",X"E6",X"E2",X"A5",X"E2",X"29",X"0F",X"C9",
		X"0A",X"B0",X"F6",X"20",X"C1",X"03",X"A5",X"E2",
		X"20",X"DC",X"FF",X"A9",X"A0",X"A8",X"20",X"EF",
		X"FF",X"A5",X"E3",X"85",X"E5",X"A5",X"E4",X"A2",
		X"05",X"94",X"E5",X"A0",X"03",X"4A",X"26",X"E5",
		X"36",X"E5",X"88",X"D0",X"F8",X"CA",X"D0",X"F1",
		X"20",X"C6",X"03",X"20",X"EF",X"FF",X"49",X"B0",
		X"C9",X"08",X"B0",X"CF",X"95",X"EF",X"CA",X"E0",
		X"FB",X"D0",X"ED",X"A0",X"FB",X"A9",X"A0",X"20",
		X"EF",X"FF",X"B5",X"F0",X"D5",X"EB",X"D0",X"0D",
		X"94",X"EB",X"A9",X"AB",X"95",X"F0",X"C8",X"D0",
		X"EE",X"A2",X"2D",X"D0",X"8B",X"E8",X"D0",X"EA",
		X"A0",X"FB",X"B6",X"F0",X"8A",X"A2",X"FB",X"D5",
		X"EB",X"D0",X"07",X"94",X"EB",X"A9",X"AD",X"20",
		X"EF",X"FF",X"E8",X"D0",X"F2",X"C8",X"D0",X"EA",
		X"F0",X"87",X"BF",X"D9",X"C4",X"C1",X"C5",X"D2",
		X"8D",X"8D",X"B7",X"AD",X"B0",X"A0",X"CD",X"CF",
		X"D2",X"C6",X"A0",X"D3",X"D4",X"C9",X"C7",X"C9",
		X"C4",X"A0",X"C5",X"D6",X"C9",X"C6",X"A0",X"D3",
		X"D3",X"C5",X"D5",X"C7",X"8D",X"8D",X"CE",X"C9",
		X"D7",X"A0",X"D5",X"CF",X"D9",X"A0",X"AB",X"A9",
		X"8D",X"4C",X"EF",X"FF",X"AD",X"11",X"D0",X"10",
		X"FB",X"AD",X"10",X"D0",X"60",X"04",X"00",X"00",
		X"D8",X"A2",X"FF",X"9A",X"A9",X"2A",X"85",X"5A",
		X"20",X"55",X"05",X"A9",X"8B",X"85",X"58",X"A9",
		X"06",X"85",X"59",X"20",X"AD",X"04",X"20",X"CB",
		X"04",X"D0",X"0E",X"A9",X"BE",X"85",X"58",X"A9",
		X"06",X"85",X"59",X"20",X"AD",X"04",X"20",X"E8",
		X"04",X"20",X"1F",X"06",X"20",X"6A",X"05",X"20",
		X"E8",X"04",X"20",X"A8",X"04",X"20",X"09",X"05",
		X"20",X"27",X"05",X"00",X"FD",X"04",X"68",X"18",
		X"20",X"BB",X"04",X"C9",X"51",X"D0",X"03",X"4C",
		X"9A",X"04",X"20",X"9E",X"05",X"A5",X"51",X"C9",
		X"10",X"D0",X"0A",X"C6",X"5D",X"F0",X"B6",X"20",
		X"38",X"05",X"4C",X"3B",X"04",X"20",X"E8",X"04",
		X"20",X"A8",X"04",X"20",X"0C",X"06",X"F0",X"03",
		X"4C",X"35",X"04",X"20",X"43",X"05",X"A9",X"8E",
		X"85",X"58",X"A9",X"07",X"85",X"59",X"20",X"AD",
		X"04",X"A5",X"55",X"20",X"EF",X"FF",X"A9",X"A3",
		X"85",X"58",X"A9",X"07",X"85",X"59",X"20",X"AD",
		X"04",X"20",X"27",X"05",X"A9",X"BB",X"85",X"58",
		X"A9",X"07",X"85",X"59",X"20",X"AD",X"04",X"20",
		X"CB",X"04",X"D0",X"03",X"4C",X"29",X"04",X"A9",
		X"D0",X"85",X"58",X"A9",X"07",X"85",X"59",X"20",
		X"AD",X"04",X"4C",X"00",X"C1",X"A9",X"0D",X"4C",
		X"EF",X"FF",X"A0",X"00",X"B1",X"58",X"F0",X"07",
		X"20",X"EF",X"FF",X"C8",X"4C",X"AF",X"04",X"60",
		X"20",X"DE",X"04",X"AD",X"11",X"D0",X"10",X"F8",
		X"AD",X"10",X"D0",X"29",X"7F",X"4C",X"EF",X"FF",
		X"20",X"BB",X"04",X"C9",X"4E",X"F0",X"0A",X"C9",
		X"59",X"F0",X"07",X"20",X"38",X"05",X"4C",X"CB",
		X"04",X"BA",X"60",X"A5",X"5A",X"0A",X"90",X"02",
		X"49",X"A9",X"85",X"5A",X"60",X"20",X"A8",X"04",
		X"20",X"A8",X"04",X"A2",X"00",X"A0",X"04",X"B5",
		X"40",X"20",X"EF",X"FF",X"88",X"D0",X"05",X"A0",
		X"04",X"20",X"A8",X"04",X"E8",X"05",X"00",X"00",
		X"E0",X"10",X"D0",X"EE",X"A9",X"08",X"85",X"5D",
		X"60",X"E6",X"56",X"A5",X"56",X"29",X"0F",X"C9",
		X"0A",X"B0",X"F6",X"A5",X"56",X"38",X"E9",X"A0",
		X"90",X"0C",X"85",X"56",X"E6",X"57",X"A5",X"57",
		X"29",X"0F",X"C9",X"0A",X"B0",X"F6",X"60",X"A5",
		X"57",X"F0",X"03",X"20",X"DC",X"FF",X"A5",X"56",
		X"20",X"DC",X"FF",X"00",X"FD",X"04",X"68",X"18",
		X"A9",X"20",X"4C",X"EF",X"FF",X"A9",X"7A",X"85",
		X"58",X"A9",X"07",X"85",X"59",X"4C",X"AD",X"04",
		X"A5",X"5A",X"29",X"38",X"AA",X"BD",X"49",X"06",
		X"F0",X"07",X"20",X"EF",X"FF",X"E8",X"4C",X"48",
		X"05",X"60",X"A9",X"20",X"85",X"4F",X"A9",X"0F",
		X"85",X"52",X"A2",X"0F",X"A0",X"4F",X"98",X"9D",
		X"3F",X"00",X"88",X"CA",X"D0",X"F8",X"60",X"A9",
		X"00",X"85",X"56",X"85",X"57",X"85",X"5C",X"A6",
		X"55",X"BD",X"13",X"06",X"85",X"5B",X"20",X"DE",
		X"04",X"A5",X"5A",X"29",X"0F",X"18",X"69",X"41",
		X"C5",X"5C",X"F0",X"F2",X"20",X"9E",X"05",X"A5",
		X"51",X"C9",X"10",X"F0",X"E9",X"A5",X"50",X"85",
		X"5C",X"C6",X"5B",X"D0",X"E1",X"20",X"0C",X"06",
		X"F0",X"CD",X"60",X"85",X"50",X"C9",X"20",X"F0",
		X"3C",X"A2",X"00",X"B5",X"40",X"C5",X"50",X"F0",
		X"08",X"E8",X"E0",X"10",X"D0",X"F5",X"4C",X"E0",
		X"05",X"86",X"51",X"8A",X"29",X"0C",X"85",X"53",
		X"A5",X"52",X"29",X"0C",X"C5",X"53",X"D0",X"10",
		X"8A",X"38",X"E5",X"52",X"10",X"05",X"A9",X"FF",
		X"4C",X"F2",X"05",X"A9",X"01",X"4C",X"F2",X"05",
		X"8A",X"29",X"03",X"85",X"53",X"A5",X"52",X"29",
		X"03",X"C5",X"53",X"F0",X"05",X"A2",X"10",X"86",
		X"51",X"60",X"8A",X"38",X"E5",X"52",X"10",X"05",
		X"A9",X"FC",X"4C",X"F2",X"05",X"A9",X"04",X"85",
		X"54",X"A5",X"52",X"AA",X"18",X"65",X"54",X"A8",
		X"B9",X"40",X"00",X"95",X"40",X"06",X"00",X"00",
		X"A9",X"20",X"99",X"40",X"00",X"84",X"52",X"C4",
		X"51",X"D0",X"E9",X"60",X"A2",X"0F",X"A9",X"4F",
		X"85",X"53",X"BD",X"3F",X"00",X"C5",X"53",X"D0",
		X"05",X"C6",X"53",X"CA",X"D0",X"F4",X"60",X"A9",
		X"60",X"85",X"58",X"A9",X"07",X"85",X"59",X"20",
		X"AD",X"04",X"20",X"00",X"FD",X"04",X"68",X"18",
		X"BB",X"04",X"85",X"55",X"C9",X"31",X"10",X"03",
		X"4C",X"3E",X"06",X"A9",X"35",X"38",X"E5",X"55",
		X"30",X"01",X"60",X"20",X"38",X"05",X"4C",X"2A",
		X"06",X"03",X"09",X"13",X"23",X"FF",X"48",X"4F",
		X"4F",X"52",X"41",X"59",X"21",X"00",X"48",X"55",
		X"5A",X"5A",X"41",X"48",X"21",X"00",X"57",X"4F",
		X"4F",X"48",X"4F",X"4F",X"21",X"00",X"59",X"49",
		X"50",X"50",X"49",X"45",X"21",X"00",X"53",X"57",
		X"45",X"45",X"54",X"21",X"00",X"00",X"43",X"4F",
		X"4F",X"4C",X"21",X"00",X"00",X"00",X"4E",X"49",
		X"43",X"45",X"21",X"00",X"00",X"00",X"47",X"41",
		X"44",X"5A",X"4F",X"4F",X"4B",X"53",X"21",X"00",
		X"0D",X"0D",X"31",X"35",X"20",X"50",X"55",X"5A",
		X"5A",X"4C",X"45",X"20",X"2D",X"20",X"42",X"59",
		X"20",X"4A",X"45",X"46",X"46",X"20",X"4A",X"45",
		X"54",X"54",X"4F",X"4E",X"0D",X"0D",X"49",X"4E",
		X"53",X"54",X"52",X"55",X"43",X"54",X"49",X"4F",
		X"4E",X"53",X"20",X"28",X"59",X"2F",X"4E",X"29",
		X"3F",X"20",X"00",X"0D",X"0D",X"54",X"59",X"50",
		X"45",X"20",X"41",X"20",X"4C",X"45",X"54",X"54",
		X"45",X"52",X"20",X"4F",X"4E",X"20",X"54",X"48",
		X"45",X"20",X"53",X"41",X"4D",X"45",X"0D",X"52",
		X"4F",X"57",X"20",X"4F",X"52",X"20",X"43",X"4F",
		X"4C",X"55",X"4D",X"4E",X"20",X"41",X"53",X"20",
		X"54",X"48",X"45",X"20",X"45",X"4D",X"50",X"54",
		X"59",X"0D",X"53",X"50",X"41",X"43",X"45",X"20",
		X"54",X"4F",X"20",X"53",X"4C",X"07",X"00",X"D8",
		X"49",X"44",X"45",X"20",X"54",X"48",X"41",X"54",
		X"20",X"4C",X"45",X"54",X"54",X"45",X"52",X"0D",
		X"28",X"41",X"4E",X"44",X"20",X"41",X"4E",X"59",
		X"20",X"42",X"45",X"54",X"57",X"45",X"45",X"4E",
		X"29",X"20",X"54",X"00",X"FD",X"04",X"68",X"18",
		X"4F",X"57",X"41",X"52",X"44",X"53",X"0D",X"54",
		X"48",X"45",X"20",X"53",X"50",X"41",X"43",X"45",
		X"2E",X"20",X"54",X"59",X"50",X"45",X"20",X"51",
		X"20",X"54",X"4F",X"20",X"51",X"55",X"49",X"54",
		X"2E",X"0D",X"54",X"48",X"49",X"53",X"20",X"49",
		X"53",X"20",X"54",X"48",X"45",X"20",X"53",X"4F",
		X"4C",X"56",X"45",X"44",X"20",X"50",X"55",X"5A",
		X"5A",X"4C",X"45",X"3A",X"00",X"0D",X"44",X"49",
		X"46",X"46",X"49",X"43",X"55",X"4C",X"54",X"59",
		X"20",X"4C",X"45",X"56",X"45",X"4C",X"20",X"28",
		X"31",X"2D",X"35",X"29",X"3F",X"20",X"00",X"0D",
		X"53",X"4F",X"52",X"52",X"59",X"2E",X"20",X"54",
		X"52",X"59",X"20",X"41",X"47",X"41",X"49",X"4E",
		X"3A",X"20",X"00",X"20",X"59",X"4F",X"55",X"20",
		X"53",X"4F",X"4C",X"56",X"45",X"44",X"0D",X"41",
		X"20",X"4C",X"45",X"56",X"45",X"4C",X"20",X"00",
		X"20",X"50",X"55",X"5A",X"5A",X"4C",X"45",X"21",
		X"0D",X"0D",X"54",X"4F",X"54",X"41",X"4C",X"20",
		X"4D",X"4F",X"56",X"45",X"53",X"3A",X"20",X"00",
		X"0D",X"0D",X"50",X"4C",X"41",X"59",X"20",X"41",
		X"47",X"41",X"49",X"4E",X"20",X"28",X"59",X"2F",
		X"4E",X"29",X"3F",X"20",X"00",X"0D",X"0D",X"42",
		X"59",X"45",X"21",X"0D",X"00",X"0B",X"E5",X"1B",
		X"20",X"EF",X"FF",X"E8",X"BD",X"F1",X"0B",X"D0",
		X"F7",X"4C",X"9D",X"0C",X"0D",X"55",X"53",X"41",
		X"47",X"45",X"3A",X"0D",X"20",X"21",X"38",X"30",
		X"30",X"3A",X"50",X"0C",X"00",X"8A",X"48",X"41",
		X"20",X"20",X"20",X"20",X"41",X"53",X"53",X"45",
		X"4D",X"42",X"4C",X"45",X"20",X"31",X"53",X"54",
		X"0D",X"20",X"21",X"20",X"4C",X"44",X"41",X"20",
		X"23",X"31",X"20",X"20",X"20",X"20",X"41",X"53",
		X"53",X"45",X"4D",X"00",X"FD",X"04",X"68",X"18",
		X"42",X"4C",X"45",X"20",X"4E",X"45",X"58",X"54",
		X"0D",X"20",X"21",X"38",X"30",X"30",X"4C",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"44",X"49",
		X"53",X"41",X"53",X"53",X"45",X"4D",X"42",X"4C",
		X"45",X"0D",X"20",X"21",X"4C",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"4E",
		X"45",X"58",X"54",X"20",X"53",X"43",X"52",X"45",
		X"45",X"4E",X"0D",X"20",X"21",X"28",X"52",X"45",
		X"54",X"55",X"52",X"4E",X"29",X"20",X"20",X"20",
		X"45",X"58",X"49",X"54",X"0D",X"20",X"42",X"45",
		X"45",X"52",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"53",X"4B",X"49",X"50",X"20",X"55",
		X"53",X"41",X"47",X"45",X"00",X"0C",X"8A",X"76",
		X"A9",X"0C",X"48",X"20",X"FD",X"0D",X"20",X"F1",
		X"0E",X"85",X"44",X"84",X"45",X"68",X"38",X"E9",
		X"01",X"D0",X"EF",X"20",X"95",X"0E",X"8A",X"D0",
		X"03",X"4C",X"1F",X"FF",X"A0",X"00",X"20",X"C0",
		X"0E",X"48",X"8A",X"F0",X"07",X"B5",X"46",X"95",
		X"44",X"CA",X"10",X"F9",X"68",X"C9",X"05",X"F0",
		X"CF",X"C9",X"99",X"F0",X"04",X"C9",X"93",X"D0",
		X"76",X"A9",X"03",X"85",X"47",X"20",X"B2",X"0E",
		X"0A",X"E9",X"BE",X"C5",X"C2",X"90",X"68",X"0A",
		X"0A",X"A2",X"04",X"0A",X"26",X"4A",X"26",X"4B",
		X"CA",X"10",X"F8",X"C6",X"47",X"F0",X"F4",X"10",
		X"E4",X"A2",X"05",X"20",X"B2",X"0E",X"84",X"3A",
		X"DD",X"52",X"0F",X"D0",X"13",X"20",X"B2",X"0E",
		X"DD",X"58",X"0F",X"F0",X"0D",X"BD",X"58",X"0F",
		X"F0",X"07",X"C9",X"A4",X"F0",X"03",X"0D",X"00",
		X"00",X"A4",X"3A",X"18",X"88",X"26",X"4C",X"E0",
		X"03",X"D0",X"0D",X"20",X"C0",X"0E",X"A5",X"49",
		X"F0",X"01",X"E8",X"86",X"38",X"A2",X"03",X"88",
		X"86",X"47",X"CA",X"00",X"FD",X"04",X"68",X"18",
		X"10",X"C9",X"A5",X"4C",X"0A",X"0A",X"05",X"38",
		X"C9",X"20",X"B0",X"06",X"A6",X"38",X"F0",X"02",
		X"09",X"80",X"85",X"4C",X"84",X"3A",X"B9",X"00",
		X"02",X"C9",X"BB",X"F0",X"04",X"C9",X"8D",X"D0",
		X"2C",X"A5",X"47",X"20",X"B7",X"0D",X"AA",X"BD",
		X"9E",X"0F",X"C5",X"4A",X"D0",X"13",X"BD",X"5E",
		X"0F",X"C5",X"4B",X"D0",X"0C",X"A5",X"4C",X"A4",
		X"40",X"C0",X"9D",X"F0",X"20",X"C5",X"40",X"F0",
		X"37",X"C6",X"47",X"D0",X"DC",X"E6",X"4C",X"C6",
		X"38",X"F0",X"D6",X"A4",X"3A",X"98",X"AA",X"20",
		X"BB",X"0E",X"20",X"79",X"0E",X"A9",X"DE",X"20",
		X"EF",X"FF",X"4C",X"9D",X"0C",X"E9",X"81",X"4A",
		X"D0",X"E9",X"A4",X"49",X"A6",X"48",X"D0",X"01",
		X"88",X"CA",X"8A",X"18",X"E5",X"44",X"85",X"48",
		X"10",X"01",X"C8",X"98",X"E5",X"45",X"D0",X"43",
		X"A4",X"41",X"B9",X"47",X"00",X"91",X"44",X"88",
		X"10",X"F8",X"A9",X"01",X"4C",X"8C",X"0C",X"A6",
		X"44",X"A4",X"45",X"20",X"BB",X"0E",X"20",X"6F",
		X"0E",X"A0",X"00",X"A9",X"AD",X"20",X"EF",X"FF",
		X"20",X"77",X"0E",X"A1",X"44",X"A8",X"4A",X"90",
		X"0B",X"4A",X"B0",X"17",X"C9",X"22",X"F0",X"13",
		X"29",X"07",X"09",X"80",X"4A",X"AA",X"BD",X"00",
		X"0F",X"B0",X"04",X"4A",X"4A",X"4A",X"4A",X"29",
		X"0F",X"D0",X"04",X"A0",X"80",X"A9",X"00",X"AA",
		X"BD",X"44",X"0F",X"85",X"40",X"29",X"03",X"85",
		X"41",X"98",X"29",X"8F",X"AA",X"98",X"A0",X"03",
		X"E0",X"8A",X"F0",X"0B",X"4A",X"90",X"08",X"4A",
		X"4A",X"09",X"20",X"88",X"D0",X"FA",X"C8",X"88",
		X"D0",X"F2",X"60",X"20",X"A1",X"0D",X"0E",X"00",
		X"00",X"48",X"B1",X"44",X"20",X"DC",X"FF",X"A2",
		X"01",X"20",X"79",X"0E",X"C4",X"41",X"C8",X"90",
		X"F1",X"A2",X"03",X"00",X"FD",X"04",X"68",X"18",
		X"C0",X"03",X"90",X"F2",X"68",X"A8",X"B9",X"5E",
		X"0F",X"85",X"42",X"B9",X"9E",X"0F",X"85",X"43",
		X"A9",X"00",X"A0",X"05",X"06",X"43",X"26",X"42",
		X"2A",X"88",X"D0",X"F8",X"69",X"BF",X"20",X"EF",
		X"FF",X"CA",X"D0",X"EC",X"20",X"77",X"0E",X"A2",
		X"06",X"E0",X"03",X"D0",X"12",X"A4",X"41",X"F0",
		X"0E",X"A5",X"40",X"C9",X"E8",X"B1",X"44",X"B0",
		X"1C",X"20",X"DC",X"FF",X"88",X"D0",X"F2",X"06",
		X"40",X"90",X"0E",X"BD",X"51",X"0F",X"20",X"EF",
		X"FF",X"BD",X"57",X"0F",X"F0",X"03",X"20",X"EF",
		X"FF",X"CA",X"D0",X"D5",X"60",X"20",X"F4",X"0E",
		X"AA",X"E8",X"D0",X"01",X"C8",X"98",X"20",X"DC",
		X"FF",X"8A",X"4C",X"DC",X"FF",X"A2",X"01",X"A9",
		X"A0",X"20",X"EF",X"FF",X"CA",X"D0",X"F8",X"60",
		X"C9",X"9B",X"F0",X"0A",X"20",X"EF",X"FF",X"C9",
		X"DF",X"F0",X"12",X"E8",X"10",X"12",X"A9",X"DC",
		X"20",X"EF",X"FF",X"20",X"BB",X"0E",X"A9",X"A1",
		X"20",X"EF",X"FF",X"A2",X"01",X"CA",X"30",X"F3",
		X"2C",X"11",X"D0",X"10",X"FB",X"AD",X"10",X"D0",
		X"9D",X"00",X"02",X"C9",X"8D",X"D0",X"D1",X"60",
		X"B9",X"00",X"02",X"C8",X"C9",X"A0",X"F0",X"F8",
		X"60",X"A9",X"8D",X"4C",X"EF",X"FF",X"A2",X"00",
		X"86",X"48",X"86",X"49",X"F0",X"15",X"A2",X"03",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"26",X"48",X"26",
		X"49",X"CA",X"10",X"F8",X"B5",X"49",X"95",X"47",
		X"E8",X"F0",X"F9",X"B9",X"00",X"02",X"C8",X"49",
		X"B0",X"C9",X"0A",X"90",X"E1",X"69",X"88",X"C9",
		X"FA",X"B0",X"DB",X"60",X"4C",X"E9",X"0B",X"A5",
		X"41",X"38",X"A4",X"45",X"AA",X"10",X"01",X"88",
		X"65",X"44",X"90",X"01",X"C8",X"60",X"0F",X"00",
		X"DE",X"40",X"02",X"45",X"03",X"D0",X"08",X"40",
		X"09",X"30",X"22",X"00",X"FD",X"04",X"68",X"18",
		X"45",X"33",X"D0",X"08",X"40",X"09",X"40",X"02",
		X"45",X"33",X"D0",X"08",X"40",X"09",X"40",X"02",
		X"45",X"B3",X"D0",X"08",X"40",X"09",X"00",X"22",
		X"44",X"33",X"D0",X"8C",X"44",X"00",X"11",X"22",
		X"44",X"33",X"D0",X"8C",X"44",X"9A",X"10",X"22",
		X"44",X"33",X"D0",X"08",X"40",X"09",X"10",X"22",
		X"44",X"33",X"D0",X"08",X"40",X"09",X"62",X"13",
		X"78",X"A9",X"00",X"21",X"81",X"82",X"00",X"00",
		X"59",X"4D",X"91",X"92",X"86",X"4A",X"85",X"9D",
		X"AC",X"A9",X"AC",X"A3",X"A8",X"A4",X"D9",X"00",
		X"D8",X"A4",X"A4",X"00",X"1C",X"8A",X"1C",X"23",
		X"5D",X"8B",X"1B",X"A1",X"9D",X"8A",X"1D",X"23",
		X"9D",X"8B",X"1D",X"A1",X"00",X"29",X"19",X"AE",
		X"69",X"A8",X"19",X"23",X"24",X"53",X"1B",X"23",
		X"24",X"53",X"19",X"A1",X"00",X"1A",X"5B",X"5B",
		X"A5",X"69",X"24",X"24",X"AE",X"AE",X"A8",X"AD",
		X"29",X"00",X"7C",X"00",X"15",X"9C",X"6D",X"9C",
		X"A5",X"69",X"29",X"53",X"84",X"13",X"34",X"11",
		X"A5",X"69",X"23",X"A0",X"D8",X"62",X"5A",X"48",
		X"26",X"62",X"94",X"88",X"54",X"44",X"C8",X"54",
		X"68",X"44",X"E8",X"94",X"00",X"B4",X"08",X"84",
		X"74",X"B4",X"28",X"6E",X"74",X"F4",X"CC",X"4A",
		X"72",X"F2",X"A4",X"8A",X"00",X"AA",X"A2",X"A2",
		X"74",X"74",X"74",X"72",X"44",X"68",X"B2",X"32",
		X"B2",X"00",X"22",X"26",X"1A",X"1A",X"26",X"26",
		X"72",X"72",X"88",X"C8",X"C4",X"CA",X"26",X"48",
		X"44",X"44",X"A2",X"C8",X"5E",X"00",X"E3",X"75",
		X"2B",X"3E",X"1A",X"3D",X"FC",X"0F",X"82",X"FF",
		X"35",X"3F",X"3B",X"11",X"10",X"D0",X"2B",X"30",
		X"1A",X"0F",X"5E",X"3D",X"8C",X"FF",X"35",X"3F",
		X"3B",X"8C",X"FF",X"E6",X"60",X"35",X"50",X"21",
		X"E6",X"20",X"E3",X"00",X"FD",X"04",X"68",X"18",
		X"60",X"8C",X"0A",X"35",X"72",X"2A",X"59",X"07",
		X"8C",X"0A",X"8C",X"1A",X"35",X"72",X"33",X"EC",
		X"00",X"8C",X"1A",X"82",X"7F",X"E6",X"80",X"F3",
		X"30",X"11",X"12",X"D0",X"2B",X"30",X"AD",X"35",
		X"3F",X"75",X"5E",X"3C",X"88",X"80",X"85",X"0F",
		X"5F",X"1A",X"1C",X"E3",X"02",X"F6",X"E3",X"42",
		X"35",X"72",X"5B",X"21",X"7A",X"E6",X"02",X"2B",
		X"7A",X"59",X"00",X"F0",X"30",X"11",X"10",X"D0",
		X"2B",X"30",X"AD",X"35",X"3F",X"6C",X"FC",X"3C",
		X"82",X"7F",X"35",X"72",X"71",X"F3",X"30",X"59",
		X"1F",X"5E",X"3C",X"1A",X"3C",X"E6",X"01",X"35",
		X"53",X"89",X"59",X"A0",X"85",X"0F",X"5F",X"21",
		X"7A",X"E6",X"06",X"2B",X"7A",X"59",X"1E",X"5E",
		X"3C",X"8C",X"14",X"35",X"72",X"9B",X"59",X"C0",
		X"85",X"0F",X"5F",X"21",X"7A",X"E6",X"06",X"2B",
		X"7A",X"11",X"07",X"5F",X"2B",X"30",X"63",X"59",
		X"FF",X"5E",X"0E",X"11",X"00",X"04",X"7F",X"3E",
		X"18",X"A2",X"00",X"A0",X"0C",X"B9",X"CE",X"5E",
		X"84",X"3A",X"A0",X"07",X"9D",X"00",X"01",X"69",
		X"01",X"E8",X"E8",X"88",X"D0",X"F6",X"E8",X"E8",
		X"E8",X"E8",X"A4",X"3A",X"88",X"10",X"E6",X"4C",
		X"05",X"C1",X"77",X"70",X"56",X"4F",X"48",X"41",
		X"3A",X"33",X"2C",X"25",X"1E",X"17",X"10",X"D8",
		X"58",X"A2",X"F7",X"9A",X"4C",X"1A",X"FF",X"5F",
		X"00",X"00",X"2B",X"1A",X"11",X"0C",X"0B",X"2B",
		X"22",X"B4",X"E6",X"11",X"FE",X"FF",X"F6",X"90",
		X"FE",X"2B",X"7C",X"DF",X"FA",X"21",X"24",X"EC",
		X"00",X"21",X"26",X"EC",X"02",X"21",X"28",X"EC",
		X"04",X"11",X"E1",X"04",X"2B",X"22",X"11",X"00",
		X"3F",X"2B",X"24",X"5E",X"26",X"21",X"7C",X"5E",
		X"27",X"8C",X"8D",X"35",X"3F",X"3B",X"1A",X"7A",
		X"E6",X"FB",X"35",X"00",X"FD",X"04",X"68",X"18",
		X"56",X"3B",X"59",X"00",X"35",X"72",X"96",X"21",
		X"7A",X"2B",X"28",X"82",X"FF",X"E6",X"FB",X"35",
		X"4D",X"4C",X"11",X"FB",X"FF",X"B4",X"CB",X"93",
		X"28",X"E3",X"01",X"35",X"50",X"4C",X"59",X"61",
		X"5E",X"7A",X"E3",X"9F",X"2B",X"7C",X"AD",X"5E",
		X"7B",X"21",X"7A",X"E6",X"02",X"2B",X"28",X"11",
		X"00",X"07",X"99",X"28",X"AD",X"82",X"01",X"5E",
		X"26",X"B4",X"CB",X"93",X"28",X"1A",X"28",X"35",
		X"72",X"66",X"21",X"7C",X"E3",X"12",X"2B",X"7E",
		X"AD",X"5E",X"26",X"21",X"7C",X"AD",X"F0",X"7E",
		X"1A",X"26",X"F0",X"7C",X"93",X"7C",X"93",X"7C",
		X"1A",X"7C",X"8C",X"D8",X"35",X"72",X"79",X"1A",
		X"27",X"E6",X"A0",X"35",X"50",X"EF",X"E6",X"40",
		X"35",X"50",X"A4",X"E6",X"20",X"E3",X"0E",X"35",
		X"53",X"B2",X"E3",X"32",X"2B",X"7C",X"11",X"00",
		X"07",X"90",X"B7",X"2B",X"7C",X"11",X"00",X"08",
		X"2B",X"7E",X"21",X"7C",X"E9",X"E9",X"99",X"7C",
		X"99",X"7E",X"2B",X"7E",X"21",X"7A",X"2B",X"28",
		X"E3",X"06",X"2B",X"7A",X"59",X"05",X"2B",X"7C",
		X"21",X"7E",X"7F",X"00",X"82",X"FE",X"5E",X"26",
		X"11",X"00",X"07",X"99",X"28",X"AD",X"35",X"3F",
		X"E2",X"93",X"26",X"B4",X"CB",X"93",X"7E",X"93",
		X"28",X"21",X"7C",X"E6",X"01",X"35",X"4D",X"CD",
		X"EE",X"00",X"2B",X"24",X"EE",X"02",X"2B",X"26",
		X"EE",X"04",X"2B",X"28",X"DF",X"06",X"FF",X"C1",
		X"00",X"58",X"A9",X"AA",X"20",X"EF",X"FF",X"AE",
		X"00",X"C2",X"BD",X"00",X"C2",X"20",X"EF",X"FF",
		X"CA",X"D0",X"F7",X"AE",X"25",X"C1",X"BD",X"25",
		X"C1",X"20",X"EF",X"FF",X"CA",X"D0",X"F7",X"2C",
		X"12",X"D0",X"30",X"FB",X"4C",X"00",X"FF",X"32",
		X"8D",X"CE",X"CF",X"CD",X"DA",X"CF",X"D7",X"A0",
		X"DA",X"AD",X"CC",X"00",X"FD",X"04",X"68",X"18",
		X"D4",X"C3",X"8D",X"D4",X"D2",X"C1",X"D4",X"D3",
		X"A0",X"CD",X"D2",X"C1",X"D7",X"A0",X"C3",X"C9",
		X"D3",X"C1",X"C2",X"A0",X"D2",X"B3",X"C2",X"B2",
		X"C5",X"8D",X"C3",X"C9",X"D3",X"C1",X"C2",X"A0",
		X"D2",X"C5",X"C7",X"C5",X"D4",X"CE",X"C9",X"C2",
		X"00",X"5B",X"5A",X"A0",X"D2",X"B0",X"B0",X"B0",
		X"C5",X"8D",X"D5",X"CE",X"C5",X"CD",X"A0",X"D2",
		X"B0",X"B0",X"B1",X"C3",X"8D",X"D2",X"C5",X"CC",
		X"C2",X"CD",X"C5",X"D3",X"D3",X"C1",X"AD",X"C9",
		X"CE",X"C9",X"CD",X"A0",X"A0",X"D2",X"C5",X"C5",
		X"C5",X"8D",X"C5",X"CC",X"DA",X"DA",X"D5",X"D0",
		X"AD",X"B5",X"B1",X"A0",X"A0",X"D2",X"B0",X"B0",
		X"B4",X"8D",X"C4",X"CE",X"C9",X"CD",X"D2",X"C5",
		X"D4",X"D3",X"C1",X"CD",X"A0",X"A0",X"D2",X"B0",
		X"B0",X"B3",X"8D",X"8D",X"CC",X"D4",X"D4",X"A0",
		X"CE",X"CF",X"A0",X"B1",X"AD",X"C5",X"CC",X"D0",
		X"D0",X"C1",X"8D",X"8D",X"8D",X"D0",X"10",X"04",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"4C",
		X"B0",X"E2",X"AD",X"11",X"D0",X"10",X"FB",X"AD",
		X"10",X"D0",X"60",X"8A",X"29",X"20",X"F0",X"23",
		X"A9",X"A0",X"85",X"44",X"4C",X"C9",X"E3",X"A9",
		X"20",X"C5",X"81",X"B0",X"0C",X"A9",X"8D",X"A0",
		X"07",X"20",X"C9",X"E3",X"A9",X"A0",X"88",X"D0",
		X"F8",X"A0",X"00",X"B1",X"42",X"E6",X"42",X"D0",
		X"02",X"E6",X"43",X"60",X"20",X"15",X"E7",X"20",
		X"76",X"E5",X"A5",X"42",X"C5",X"46",X"A5",X"43",
		X"E5",X"47",X"B0",X"EF",X"20",X"6D",X"E0",X"4C",
		X"3B",X"E0",X"A5",X"CA",X"85",X"42",X"A5",X"CB",
		X"85",X"43",X"A5",X"4C",X"85",X"46",X"A5",X"4D",
		X"85",X"47",X"D0",X"DE",X"20",X"15",X"E7",X"20",
		X"6D",X"E5",X"A5",X"44",X"85",X"42",X"A5",X"45",
		X"85",X"43",X"B0",X"00",X"FD",X"04",X"68",X"18",
		X"C7",X"86",X"D8",X"A9",X"A0",X"85",X"82",X"20",
		X"2A",X"E0",X"98",X"85",X"44",X"20",X"2A",X"E0",
		X"AA",X"20",X"2A",X"E0",X"20",X"1B",X"E5",X"20",
		X"18",X"E0",X"84",X"82",X"AA",X"10",X"18",X"0A",
		X"10",X"E9",X"A5",X"44",X"D0",X"03",X"20",X"11",
		X"E0",X"8A",X"20",X"C9",X"E3",X"A9",X"25",X"20",
		X"1A",X"E0",X"AA",X"30",X"F5",X"85",X"44",X"C9",
		X"01",X"D0",X"05",X"A6",X"D8",X"4C",X"CD",X"E3",
		X"48",X"84",X"CE",X"A2",X"ED",X"86",X"CF",X"C9",
		X"51",X"90",X"04",X"C6",X"CF",X"E9",X"50",X"48",
		X"B1",X"CE",X"AA",X"88",X"B1",X"CE",X"10",X"FA",
		X"E0",X"C0",X"B0",X"04",X"E0",X"00",X"30",X"F2",
		X"AA",X"68",X"E9",X"01",X"D0",X"E9",X"24",X"44",
		X"30",X"03",X"20",X"F8",X"EF",X"B1",X"CE",X"10",
		X"10",X"AA",X"29",X"3F",X"85",X"44",X"18",X"69",
		X"A0",X"20",X"C9",X"E3",X"88",X"E0",X"C0",X"90",
		X"EC",X"20",X"0C",X"E0",X"68",X"C9",X"5D",X"F0",
		X"A4",X"C9",X"28",X"D0",X"8A",X"F0",X"9E",X"20",
		X"18",X"E1",X"95",X"50",X"E1",X"00",X"00",X"D5",
		X"88",X"90",X"11",X"A0",X"2B",X"4C",X"E0",X"E3",
		X"20",X"34",X"EE",X"D5",X"50",X"90",X"F4",X"20",
		X"E4",X"EF",X"95",X"88",X"4C",X"23",X"E8",X"20",
		X"34",X"EE",X"F0",X"E7",X"38",X"E9",X"01",X"60",
		X"20",X"18",X"E1",X"95",X"50",X"18",X"F5",X"88",
		X"4C",X"02",X"E1",X"A0",X"14",X"D0",X"D6",X"20",
		X"18",X"E1",X"E8",X"B5",X"50",X"85",X"DA",X"65",
		X"CE",X"48",X"A8",X"B5",X"88",X"85",X"DB",X"65",
		X"CF",X"48",X"C4",X"CA",X"E5",X"CB",X"B0",X"E3",
		X"A5",X"DA",X"69",X"FE",X"85",X"DA",X"A9",X"FF",
		X"A8",X"65",X"DB",X"85",X"DB",X"C8",X"B1",X"DA",
		X"D9",X"CC",X"00",X"D0",X"0F",X"98",X"F0",X"F5",
		X"68",X"91",X"DA",X"00",X"FD",X"04",X"68",X"18",
		X"99",X"CC",X"00",X"88",X"10",X"F7",X"E8",X"60",
		X"EA",X"A0",X"80",X"D0",X"95",X"A9",X"00",X"20",
		X"0A",X"E7",X"A0",X"02",X"94",X"88",X"20",X"0A",
		X"E7",X"A9",X"BF",X"20",X"C9",X"E3",X"A0",X"00",
		X"20",X"9E",X"E2",X"94",X"88",X"EA",X"EA",X"EA",
		X"B5",X"51",X"85",X"CE",X"B5",X"89",X"85",X"CF",
		X"E8",X"E8",X"20",X"BC",X"E1",X"B5",X"4E",X"D5",
		X"86",X"B0",X"15",X"F6",X"4E",X"A8",X"B1",X"CE",
		X"B4",X"50",X"C4",X"44",X"90",X"04",X"A0",X"83",
		X"D0",X"C1",X"91",X"DA",X"F6",X"50",X"90",X"E5",
		X"B4",X"50",X"8A",X"91",X"DA",X"E8",X"E8",X"60",
		X"B5",X"51",X"85",X"DA",X"38",X"E9",X"02",X"85",
		X"44",X"B5",X"89",X"85",X"DB",X"E9",X"00",X"85",
		X"45",X"A0",X"00",X"B1",X"44",X"18",X"E5",X"DA",
		X"85",X"44",X"60",X"B5",X"53",X"85",X"CE",X"B5",
		X"8B",X"85",X"CF",X"B5",X"51",X"85",X"DA",X"B5",
		X"89",X"85",X"DB",X"E8",X"E8",X"E8",X"A0",X"00",
		X"94",X"88",X"94",X"A8",X"C8",X"94",X"50",X"B5",
		X"4D",X"D5",X"85",X"08",X"48",X"B5",X"4F",X"D5",
		X"87",X"90",X"07",X"68",X"E2",X"00",X"00",X"28",
		X"B0",X"02",X"56",X"50",X"60",X"A8",X"B1",X"CE",
		X"85",X"44",X"68",X"A8",X"28",X"B0",X"F3",X"B1",
		X"DA",X"C5",X"44",X"D0",X"ED",X"F6",X"4F",X"F6",
		X"4D",X"B0",X"D7",X"20",X"D7",X"E1",X"4C",X"36",
		X"E7",X"20",X"54",X"E2",X"06",X"CE",X"26",X"CF",
		X"90",X"0D",X"18",X"A5",X"46",X"65",X"DA",X"85",
		X"46",X"A5",X"47",X"65",X"DB",X"85",X"47",X"88",
		X"F0",X"09",X"06",X"46",X"26",X"47",X"10",X"E4",
		X"4C",X"7E",X"E7",X"A5",X"46",X"20",X"08",X"E7",
		X"A5",X"47",X"95",X"A8",X"06",X"45",X"90",X"28",
		X"4C",X"6F",X"E7",X"A9",X"55",X"85",X"45",X"20",
		X"5B",X"E2",X"A5",X"00",X"FD",X"04",X"68",X"18",
		X"CE",X"85",X"DA",X"A5",X"CF",X"85",X"DB",X"20",
		X"15",X"E7",X"84",X"46",X"84",X"47",X"A5",X"CF",
		X"10",X"09",X"CA",X"06",X"45",X"20",X"6F",X"E7",
		X"20",X"15",X"E7",X"A0",X"10",X"60",X"20",X"6C",
		X"EE",X"F0",X"C5",X"FF",X"C9",X"84",X"D0",X"02",
		X"46",X"78",X"C9",X"DF",X"F0",X"11",X"C9",X"9B",
		X"F0",X"06",X"99",X"00",X"02",X"C8",X"10",X"0A",
		X"A0",X"8B",X"20",X"C4",X"E3",X"A0",X"01",X"88",
		X"30",X"F6",X"20",X"03",X"E0",X"EA",X"EA",X"20",
		X"C9",X"E3",X"C9",X"8D",X"D0",X"D6",X"A9",X"DF",
		X"99",X"00",X"02",X"60",X"20",X"D3",X"EF",X"20",
		X"CD",X"E3",X"46",X"D9",X"A9",X"BE",X"20",X"C9",
		X"E3",X"A0",X"00",X"84",X"82",X"24",X"78",X"10",
		X"0C",X"A6",X"76",X"A5",X"77",X"20",X"1B",X"E5",
		X"A9",X"A0",X"20",X"C9",X"E3",X"A2",X"FF",X"9A",
		X"20",X"9E",X"E2",X"84",X"E9",X"8A",X"85",X"C8",
		X"A2",X"18",X"20",X"91",X"E4",X"A5",X"C8",X"69",
		X"00",X"85",X"DE",X"A9",X"00",X"AA",X"69",X"02",
		X"85",X"DF",X"A1",X"DE",X"29",X"F0",X"C9",X"B0",
		X"F0",X"03",X"4C",X"83",X"E8",X"A0",X"02",X"B1",
		X"DE",X"99",X"CD",X"00",X"E3",X"00",X"00",X"88",
		X"D0",X"F8",X"20",X"8A",X"E3",X"A5",X"E9",X"E5",
		X"C8",X"C9",X"04",X"F0",X"A8",X"91",X"DE",X"A5",
		X"CA",X"F1",X"DE",X"85",X"44",X"A5",X"CB",X"E9",
		X"00",X"85",X"45",X"A5",X"44",X"C5",X"CC",X"A5",
		X"45",X"E5",X"CD",X"90",X"45",X"A5",X"CA",X"F1",
		X"DE",X"85",X"46",X"A5",X"CB",X"E9",X"00",X"85",
		X"47",X"B1",X"CA",X"91",X"46",X"E6",X"CA",X"D0",
		X"02",X"E6",X"CB",X"A5",X"42",X"C5",X"CA",X"A5",
		X"43",X"E5",X"CB",X"B0",X"E0",X"B5",X"44",X"95",
		X"CA",X"CA",X"10",X"F9",X"B1",X"DE",X"A8",X"88",
		X"B1",X"DE",X"91",X"00",X"FD",X"04",X"68",X"18",
		X"46",X"98",X"D0",X"F8",X"24",X"78",X"10",X"09",
		X"B5",X"77",X"75",X"75",X"95",X"77",X"E8",X"F0",
		X"F7",X"10",X"7E",X"00",X"00",X"00",X"00",X"A0",
		X"14",X"D0",X"71",X"20",X"15",X"E7",X"A5",X"42",
		X"85",X"46",X"A5",X"43",X"85",X"47",X"20",X"75",
		X"E5",X"A5",X"42",X"85",X"44",X"A5",X"43",X"85",
		X"45",X"D0",X"0E",X"20",X"15",X"E7",X"20",X"6D",
		X"E5",X"A5",X"46",X"85",X"42",X"A5",X"47",X"85",
		X"43",X"A0",X"00",X"A5",X"CA",X"C5",X"44",X"A5",
		X"CB",X"E5",X"45",X"B0",X"16",X"A5",X"44",X"D0",
		X"02",X"C6",X"45",X"C6",X"44",X"A5",X"46",X"D0",
		X"02",X"C6",X"47",X"C6",X"46",X"B1",X"44",X"91",
		X"46",X"90",X"E0",X"A5",X"46",X"85",X"CA",X"A5",
		X"47",X"85",X"CB",X"60",X"20",X"C9",X"E3",X"C8",
		X"B9",X"00",X"EB",X"30",X"F7",X"C9",X"8D",X"D0",
		X"06",X"A9",X"00",X"85",X"81",X"A9",X"8D",X"E6",
		X"81",X"4C",X"EF",X"FF",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"A0",X"06",X"20",X"D3",X"EE",X"24",
		X"D9",X"30",X"03",X"4C",X"B6",X"E2",X"4C",X"9A",
		X"EB",X"2A",X"69",X"A0",X"DD",X"00",X"02",X"D0",
		X"53",X"B1",X"86",X"0A",X"30",X"06",X"88",X"B1",
		X"86",X"30",X"29",X"C8",X"E4",X"00",X"00",X"86",
		X"C8",X"98",X"48",X"A2",X"00",X"A1",X"86",X"AA",
		X"4A",X"49",X"48",X"11",X"86",X"C9",X"C0",X"90",
		X"01",X"E8",X"C8",X"D0",X"F3",X"68",X"A8",X"8A",
		X"4C",X"C0",X"E4",X"E6",X"E9",X"A6",X"E9",X"F0",
		X"BC",X"9D",X"00",X"02",X"60",X"A6",X"C8",X"A9",
		X"A0",X"E8",X"DD",X"00",X"02",X"B0",X"FA",X"B1",
		X"86",X"29",X"3F",X"4A",X"D0",X"B6",X"BD",X"00",
		X"02",X"B0",X"06",X"69",X"3F",X"C9",X"1A",X"90",
		X"6F",X"69",X"4F",X"C9",X"0A",X"90",X"69",X"A6",
		X"85",X"C8",X"B1",X"00",X"FD",X"04",X"68",X"18",
		X"86",X"29",X"E0",X"C9",X"20",X"F0",X"7A",X"B5",
		X"B0",X"85",X"C8",X"B5",X"D1",X"85",X"E9",X"88",
		X"B1",X"86",X"0A",X"10",X"FA",X"88",X"B0",X"38",
		X"0A",X"30",X"35",X"B4",X"58",X"84",X"87",X"B4",
		X"90",X"E8",X"10",X"DA",X"F0",X"B3",X"C9",X"7E",
		X"B0",X"22",X"CA",X"10",X"04",X"A0",X"06",X"10",
		X"29",X"94",X"90",X"A4",X"87",X"94",X"58",X"A4",
		X"C8",X"94",X"B0",X"A4",X"E9",X"94",X"D1",X"29",
		X"1F",X"A8",X"B9",X"20",X"EC",X"0A",X"A8",X"A9",
		X"76",X"2A",X"85",X"87",X"D0",X"01",X"C8",X"C8",
		X"86",X"85",X"B1",X"86",X"30",X"84",X"D0",X"05",
		X"A0",X"0E",X"4C",X"E0",X"E3",X"C9",X"03",X"B0",
		X"C3",X"4A",X"A6",X"C8",X"E8",X"BD",X"00",X"02",
		X"90",X"04",X"C9",X"A2",X"F0",X"0A",X"C9",X"DF",
		X"F0",X"06",X"86",X"C8",X"20",X"1C",X"E4",X"C8",
		X"88",X"A6",X"85",X"B1",X"86",X"88",X"0A",X"10",
		X"CF",X"B4",X"58",X"84",X"87",X"B4",X"90",X"E8",
		X"B1",X"86",X"29",X"9F",X"D0",X"ED",X"85",X"72",
		X"85",X"73",X"98",X"48",X"86",X"85",X"B4",X"D0",
		X"84",X"C9",X"18",X"A9",X"0A",X"85",X"79",X"A2",
		X"00",X"C8",X"B9",X"00",X"02",X"29",X"0F",X"65",
		X"72",X"48",X"8A",X"65",X"73",X"30",X"1C",X"AA",
		X"68",X"C6",X"79",X"D0",X"E5",X"00",X"00",X"F2",
		X"85",X"72",X"86",X"73",X"C4",X"E9",X"D0",X"DE",
		X"A4",X"C9",X"C8",X"84",X"E9",X"20",X"1C",X"E4",
		X"68",X"A8",X"A5",X"73",X"B0",X"A9",X"A0",X"00",
		X"10",X"8B",X"85",X"73",X"86",X"72",X"A2",X"04",
		X"86",X"C9",X"A9",X"B0",X"85",X"79",X"A5",X"72",
		X"DD",X"63",X"E5",X"A5",X"73",X"FD",X"68",X"E5",
		X"90",X"0D",X"85",X"73",X"A5",X"72",X"FD",X"63",
		X"E5",X"85",X"72",X"E6",X"79",X"D0",X"E7",X"A5",
		X"79",X"E8",X"CA",X"00",X"FD",X"04",X"68",X"18",
		X"F0",X"0E",X"C9",X"B0",X"F0",X"02",X"85",X"C9",
		X"24",X"C9",X"30",X"04",X"A5",X"82",X"F0",X"0B",
		X"20",X"C9",X"E3",X"24",X"78",X"10",X"04",X"99",
		X"00",X"02",X"C8",X"CA",X"10",X"C1",X"60",X"01",
		X"0A",X"64",X"E8",X"10",X"00",X"00",X"00",X"03",
		X"27",X"A5",X"CA",X"85",X"46",X"A5",X"CB",X"85",
		X"47",X"E8",X"A5",X"47",X"85",X"45",X"A5",X"46",
		X"85",X"44",X"C5",X"4C",X"A5",X"45",X"E5",X"4D",
		X"B0",X"26",X"A0",X"01",X"B1",X"44",X"E5",X"CE",
		X"C8",X"B1",X"44",X"E5",X"CF",X"B0",X"19",X"A0",
		X"00",X"A5",X"46",X"71",X"44",X"85",X"46",X"90",
		X"03",X"E6",X"47",X"18",X"C8",X"A5",X"CE",X"F1",
		X"44",X"C8",X"A5",X"CF",X"F1",X"44",X"B0",X"CA",
		X"60",X"46",X"78",X"A5",X"4C",X"85",X"CA",X"A5",
		X"4D",X"85",X"CB",X"A5",X"4A",X"85",X"CC",X"A5",
		X"4B",X"85",X"CD",X"A9",X"00",X"85",X"83",X"85",
		X"84",X"85",X"86",X"A9",X"00",X"85",X"1D",X"60",
		X"A5",X"D0",X"69",X"05",X"85",X"D2",X"A5",X"D1",
		X"69",X"00",X"85",X"D3",X"A5",X"D2",X"C5",X"CA",
		X"A5",X"D3",X"E5",X"CB",X"90",X"03",X"4C",X"6B",
		X"E3",X"A5",X"CE",X"91",X"D0",X"A5",X"CF",X"C8",
		X"91",X"D0",X"A5",X"D2",X"C8",X"91",X"D0",X"A5",
		X"D3",X"C8",X"91",X"D0",X"A9",X"00",X"C8",X"91",
		X"D0",X"C8",X"91",X"D0",X"E6",X"00",X"00",X"A5",
		X"D2",X"85",X"CC",X"A5",X"D3",X"85",X"CD",X"A5",
		X"D0",X"90",X"43",X"85",X"CE",X"84",X"CF",X"20",
		X"FF",X"E6",X"30",X"0E",X"C9",X"40",X"F0",X"0A",
		X"4C",X"28",X"E6",X"06",X"C9",X"49",X"D0",X"07",
		X"A9",X"49",X"85",X"CF",X"20",X"FF",X"E6",X"A5",
		X"4B",X"85",X"D1",X"A5",X"4A",X"85",X"D0",X"C5",
		X"CC",X"A5",X"D1",X"E5",X"CD",X"B0",X"94",X"B1",
		X"D0",X"C8",X"C5",X"00",X"FD",X"04",X"68",X"18",
		X"CE",X"D0",X"06",X"B1",X"D0",X"C5",X"CF",X"F0",
		X"0E",X"C8",X"B1",X"D0",X"48",X"C8",X"B1",X"D0",
		X"85",X"D1",X"68",X"A0",X"00",X"F0",X"DB",X"A5",
		X"D0",X"69",X"03",X"20",X"0A",X"E7",X"A5",X"D1",
		X"69",X"00",X"95",X"88",X"A5",X"CF",X"C9",X"40",
		X"D0",X"1C",X"88",X"98",X"20",X"0A",X"E7",X"88",
		X"94",X"88",X"A0",X"03",X"F6",X"88",X"C8",X"B1",
		X"D0",X"30",X"F9",X"10",X"09",X"A9",X"00",X"85",
		X"D4",X"85",X"D5",X"A2",X"18",X"48",X"A0",X"00",
		X"B1",X"DE",X"10",X"18",X"0A",X"30",X"81",X"20",
		X"FF",X"E6",X"20",X"08",X"E7",X"20",X"FF",X"E6",
		X"95",X"A8",X"24",X"D4",X"10",X"01",X"CA",X"20",
		X"FF",X"E6",X"B0",X"E6",X"C9",X"28",X"D0",X"1F",
		X"A5",X"DE",X"20",X"0A",X"E7",X"A5",X"DF",X"95",
		X"88",X"24",X"D4",X"30",X"0B",X"A9",X"01",X"20",
		X"0A",X"E7",X"A9",X"00",X"95",X"88",X"F6",X"88",
		X"20",X"FF",X"E6",X"30",X"F9",X"B0",X"D3",X"24",
		X"D4",X"10",X"06",X"C9",X"04",X"B0",X"D0",X"46",
		X"D4",X"A8",X"85",X"D6",X"B9",X"98",X"E9",X"29",
		X"55",X"0A",X"85",X"D7",X"68",X"A8",X"B9",X"98",
		X"E9",X"29",X"AA",X"C5",X"D7",X"B0",X"09",X"98",
		X"48",X"20",X"FF",X"E6",X"A5",X"D6",X"90",X"95",
		X"B9",X"10",X"EA",X"85",X"CE",X"B9",X"88",X"EA",
		X"85",X"CF",X"20",X"FC",X"E6",X"4C",X"D8",X"E6",
		X"6C",X"CE",X"00",X"E6",X"E7",X"00",X"00",X"DE",
		X"D0",X"02",X"E6",X"DF",X"B1",X"DE",X"60",X"94",
		X"87",X"CA",X"30",X"03",X"95",X"50",X"60",X"A0",
		X"66",X"4C",X"E0",X"E3",X"A0",X"00",X"B5",X"50",
		X"85",X"CE",X"B5",X"A8",X"85",X"CF",X"B5",X"88",
		X"F0",X"0E",X"85",X"CF",X"B1",X"CE",X"48",X"C8",
		X"B1",X"CE",X"85",X"CF",X"68",X"85",X"CE",X"88",
		X"E8",X"60",X"20",X"00",X"FD",X"04",X"68",X"18",
		X"4A",X"E7",X"20",X"15",X"E7",X"98",X"20",X"08",
		X"E7",X"95",X"A8",X"C5",X"CE",X"D0",X"06",X"C5",
		X"CF",X"D0",X"02",X"F6",X"50",X"60",X"20",X"82",
		X"E7",X"20",X"59",X"E7",X"20",X"15",X"E7",X"24",
		X"CF",X"30",X"1B",X"CA",X"60",X"20",X"15",X"E7",
		X"A5",X"CF",X"D0",X"04",X"A5",X"CE",X"F0",X"F3",
		X"A9",X"FF",X"20",X"08",X"E7",X"95",X"A8",X"24",
		X"CF",X"30",X"E9",X"20",X"15",X"E7",X"98",X"38",
		X"E5",X"CE",X"20",X"08",X"E7",X"98",X"E5",X"CF",
		X"50",X"23",X"A0",X"00",X"10",X"90",X"20",X"6F",
		X"E7",X"20",X"15",X"E7",X"A5",X"CE",X"85",X"DA",
		X"A5",X"CF",X"85",X"DB",X"20",X"15",X"E7",X"18",
		X"A5",X"CE",X"65",X"DA",X"20",X"08",X"E7",X"A5",
		X"CF",X"65",X"DB",X"70",X"DD",X"95",X"A8",X"60",
		X"20",X"15",X"E7",X"A4",X"CE",X"F0",X"05",X"88",
		X"A5",X"CF",X"F0",X"0C",X"60",X"A5",X"81",X"09",
		X"07",X"A8",X"C8",X"A9",X"A0",X"20",X"C9",X"E3",
		X"C4",X"81",X"B0",X"F7",X"60",X"20",X"B1",X"E7",
		X"20",X"15",X"E7",X"A5",X"CF",X"10",X"0A",X"A9",
		X"AD",X"20",X"C9",X"E3",X"20",X"72",X"E7",X"50",
		X"EF",X"88",X"84",X"D5",X"86",X"CF",X"A6",X"CE",
		X"20",X"1B",X"E5",X"A6",X"CF",X"60",X"20",X"15",
		X"E7",X"A5",X"CE",X"85",X"76",X"A5",X"CF",X"85",
		X"77",X"88",X"84",X"78",X"C8",X"A9",X"0A",X"85",
		X"74",X"84",X"75",X"60",X"20",X"15",X"E7",X"A5",
		X"CE",X"A4",X"CF",X"10",X"E8",X"00",X"00",X"F2",
		X"20",X"15",X"E7",X"B5",X"50",X"85",X"DA",X"B5",
		X"88",X"85",X"DB",X"A5",X"CE",X"91",X"DA",X"C8",
		X"A5",X"CF",X"91",X"DA",X"E8",X"60",X"68",X"68",
		X"24",X"D5",X"10",X"05",X"20",X"CD",X"E3",X"46",
		X"D5",X"60",X"A0",X"FF",X"84",X"D7",X"60",X"20",
		X"CD",X"EF",X"F0",X"00",X"FD",X"04",X"68",X"18",
		X"07",X"A9",X"25",X"85",X"D6",X"88",X"84",X"D4",
		X"E8",X"60",X"A5",X"CA",X"A4",X"CB",X"D0",X"5A",
		X"A0",X"41",X"A5",X"84",X"C9",X"08",X"B0",X"5E",
		X"A8",X"E6",X"84",X"A5",X"DE",X"99",X"00",X"11",
		X"A5",X"DF",X"99",X"08",X"11",X"A5",X"DC",X"99",
		X"10",X"11",X"A5",X"DD",X"99",X"18",X"11",X"20",
		X"15",X"E7",X"20",X"6D",X"E5",X"90",X"04",X"A0",
		X"37",X"D0",X"3B",X"A5",X"44",X"A4",X"45",X"85",
		X"DC",X"84",X"DD",X"2C",X"11",X"D0",X"30",X"4F",
		X"18",X"69",X"03",X"90",X"01",X"C8",X"A2",X"FF",
		X"86",X"D9",X"9A",X"85",X"DE",X"84",X"DF",X"20",
		X"79",X"E6",X"24",X"D9",X"10",X"49",X"18",X"A0",
		X"00",X"A5",X"DC",X"71",X"DC",X"A4",X"DD",X"90",
		X"01",X"C8",X"C5",X"4C",X"D0",X"D1",X"C4",X"4D",
		X"D0",X"CD",X"A0",X"34",X"46",X"D9",X"4C",X"E0",
		X"E3",X"A0",X"4A",X"A5",X"84",X"F0",X"F7",X"C6",
		X"84",X"A8",X"B9",X"0F",X"11",X"85",X"DC",X"B9",
		X"17",X"11",X"85",X"DD",X"BE",X"87",X"00",X"B9",
		X"07",X"11",X"A8",X"8A",X"4C",X"7A",X"E8",X"A0",
		X"63",X"20",X"C4",X"E3",X"A0",X"01",X"B1",X"DC",
		X"AA",X"C8",X"B1",X"DC",X"20",X"1B",X"E5",X"4C",
		X"B3",X"E2",X"C6",X"83",X"A0",X"5B",X"A5",X"83",
		X"F0",X"C4",X"A8",X"B5",X"50",X"D9",X"FF",X"11",
		X"D0",X"F0",X"B5",X"88",X"D9",X"07",X"12",X"D0",
		X"E9",X"B9",X"0F",X"12",X"85",X"DA",X"B9",X"17",
		X"12",X"85",X"DB",X"20",X"15",X"E7",X"CA",X"20",
		X"93",X"E7",X"20",X"01",X"E9",X"00",X"00",X"E8",
		X"CA",X"A4",X"83",X"B9",X"47",X"12",X"95",X"A7",
		X"B9",X"3F",X"12",X"A0",X"00",X"20",X"08",X"E7",
		X"20",X"82",X"E7",X"20",X"59",X"E7",X"20",X"15",
		X"E7",X"A4",X"83",X"A5",X"CE",X"F0",X"05",X"59",
		X"17",X"12",X"10",X"00",X"FD",X"04",X"68",X"18",
		X"12",X"B9",X"1F",X"12",X"85",X"DC",X"B9",X"27",
		X"12",X"85",X"DD",X"BE",X"2F",X"12",X"B9",X"37",
		X"12",X"D0",X"87",X"C6",X"83",X"60",X"A0",X"54",
		X"A5",X"83",X"C9",X"08",X"F0",X"9A",X"E6",X"83",
		X"A8",X"B5",X"50",X"99",X"00",X"12",X"B5",X"88",
		X"99",X"08",X"12",X"60",X"20",X"15",X"E7",X"A4",
		X"83",X"A5",X"CE",X"99",X"3F",X"12",X"A5",X"CF",
		X"99",X"47",X"12",X"A9",X"01",X"99",X"0F",X"12",
		X"A9",X"00",X"99",X"17",X"12",X"A5",X"DC",X"99",
		X"1F",X"12",X"A5",X"DD",X"99",X"27",X"12",X"A5",
		X"DE",X"99",X"2F",X"12",X"A5",X"DF",X"99",X"37",
		X"12",X"60",X"20",X"15",X"E7",X"A4",X"83",X"A5",
		X"CE",X"99",X"0F",X"12",X"A5",X"CF",X"4C",X"66",
		X"E9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"3F",X"3F",
		X"C0",X"C0",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",
		X"3C",X"30",X"0F",X"C0",X"CC",X"FF",X"55",X"00",
		X"AB",X"AB",X"03",X"03",X"FF",X"FF",X"55",X"FF",
		X"FF",X"55",X"CF",X"CF",X"CF",X"CF",X"CF",X"FF",
		X"55",X"C3",X"C3",X"C3",X"55",X"F0",X"F0",X"CF",
		X"56",X"56",X"56",X"55",X"FF",X"FF",X"55",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"00",X"AB",X"03",X"57",X"03",X"03",X"03",
		X"03",X"07",X"03",X"03",X"EA",X"00",X"00",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",
		X"03",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"17",
		X"FF",X"FF",X"19",X"5D",X"35",X"4B",X"F2",X"EC",
		X"87",X"6F",X"AD",X"00",X"FD",X"04",X"68",X"18",
		X"B7",X"E2",X"F8",X"54",X"80",X"96",X"85",X"82",
		X"22",X"10",X"33",X"4A",X"13",X"06",X"0B",X"4A",
		X"01",X"40",X"47",X"7A",X"00",X"FF",X"23",X"09",
		X"5B",X"16",X"B6",X"CB",X"FF",X"FF",X"FB",X"FF",
		X"FF",X"24",X"F6",X"4E",X"59",X"50",X"00",X"FF",
		X"23",X"A3",X"6F",X"36",X"23",X"D7",X"1C",X"22",
		X"C2",X"AE",X"BA",X"23",X"FF",X"FF",X"21",X"30",
		X"1E",X"03",X"C4",X"20",X"00",X"C1",X"FF",X"FF",
		X"FF",X"A0",X"30",X"1E",X"A4",X"D3",X"B6",X"BC",
		X"AA",X"3A",X"01",X"50",X"7E",X"D8",X"D8",X"A5",
		X"3C",X"FF",X"16",X"5B",X"28",X"03",X"C4",X"1D",
		X"00",X"0C",X"4E",X"00",X"3E",X"00",X"A6",X"B0",
		X"00",X"BC",X"C6",X"57",X"8C",X"01",X"27",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"E8",X"FF",X"FF",X"E8",
		X"E0",X"E0",X"E0",X"EF",X"EF",X"E3",X"E3",X"E5",
		X"E5",X"E7",X"E7",X"EE",X"EF",X"EF",X"E7",X"E7",
		X"E2",X"EF",X"E7",X"E7",X"EC",X"EC",X"EC",X"E7",
		X"EC",X"EC",X"EC",X"E2",X"00",X"FF",X"E8",X"E1",
		X"E8",X"E8",X"EF",X"EB",X"FF",X"FF",X"E0",X"FF",
		X"FF",X"EF",X"EE",X"EF",X"E7",X"E7",X"00",X"FF",
		X"E8",X"E7",X"E7",X"E7",X"E8",X"E1",X"E2",X"EE",
		X"EE",X"EE",X"EE",X"E8",X"FF",X"FF",X"E1",X"E1",
		X"EF",X"EE",X"E7",X"E8",X"EE",X"E7",X"FF",X"FF",
		X"FF",X"EE",X"E1",X"EF",X"E7",X"E8",X"EF",X"EF",
		X"EB",X"E9",X"E8",X"E9",X"E9",X"E8",X"E8",X"E8",
		X"E8",X"FF",X"E8",X"E8",X"E8",X"EE",X"E7",X"E8",
		X"EF",X"EF",X"EE",X"EF",X"EE",X"EF",X"EE",X"EE",
		X"EF",X"EE",X"EE",X"EE",X"E1",X"E8",X"E8",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"EB",X"00",X"00",X"BE",
		X"B3",X"B2",X"B7",X"B6",X"37",X"D4",X"CF",X"CF",
		X"A0",X"CC",X"CF",X"CE",X"47",X"D3",X"D9",X"CE",
		X"D4",X"C1",X"58",X"00",X"FD",X"04",X"68",X"18",
		X"CD",X"C5",X"CD",X"A0",X"C6",X"D5",X"CC",X"4C",
		X"D4",X"CF",X"CF",X"A0",X"CD",X"C1",X"CE",X"D9",
		X"A0",X"D0",X"C1",X"D2",X"C5",X"CE",X"53",X"D3",
		X"D4",X"D2",X"C9",X"CE",X"47",X"CE",X"CF",X"A0",
		X"C5",X"CE",X"44",X"C2",X"C1",X"C4",X"A0",X"C2",
		X"D2",X"C1",X"CE",X"C3",X"48",X"BE",X"B8",X"A0",
		X"C7",X"CF",X"D3",X"D5",X"C2",X"53",X"C2",X"C1",
		X"C4",X"A0",X"D2",X"C5",X"D4",X"D5",X"D2",X"4E",
		X"BE",X"B8",X"A0",X"C6",X"CF",X"D2",X"53",X"C2",
		X"C1",X"C4",X"A0",X"CE",X"C5",X"D8",X"54",X"D3",
		X"D4",X"CF",X"D0",X"D0",X"C5",X"C4",X"A0",X"C1",
		X"D4",X"20",X"AA",X"AA",X"AA",X"20",X"A0",X"C5",
		X"D2",X"D2",X"0D",X"BE",X"B2",X"B5",X"35",X"D2",
		X"C1",X"CE",X"C7",X"45",X"C4",X"C9",X"4D",X"D3",
		X"D4",X"D2",X"A0",X"CF",X"D6",X"C6",X"4C",X"DC",
		X"0D",X"D2",X"C5",X"D4",X"D9",X"D0",X"C5",X"A0",
		X"CC",X"C9",X"CE",X"C5",X"8D",X"3F",X"46",X"D9",
		X"90",X"03",X"4C",X"C3",X"E8",X"A6",X"CF",X"9A",
		X"A6",X"CE",X"A0",X"8D",X"D0",X"02",X"A0",X"99",
		X"20",X"C4",X"E3",X"86",X"CE",X"BA",X"86",X"CF",
		X"A0",X"FE",X"84",X"D9",X"C8",X"84",X"C8",X"20",
		X"99",X"E2",X"84",X"E9",X"A2",X"18",X"A9",X"30",
		X"20",X"91",X"E4",X"E6",X"D9",X"A6",X"CE",X"A4",
		X"C8",X"0A",X"85",X"CE",X"C8",X"B9",X"00",X"02",
		X"C9",X"74",X"F0",X"D2",X"49",X"B0",X"C9",X"0A",
		X"B0",X"F0",X"C8",X"C8",X"84",X"C8",X"B9",X"00",
		X"02",X"48",X"B9",X"FF",X"01",X"A0",X"00",X"20",
		X"08",X"E7",X"68",X"95",X"A8",X"A5",X"CE",X"C9",
		X"C7",X"D0",X"03",X"20",X"6F",X"E7",X"4C",X"01",
		X"E8",X"FF",X"FF",X"FF",X"EC",X"00",X"00",X"50",
		X"20",X"13",X"EC",X"D0",X"15",X"20",X"0B",X"EC",
		X"D0",X"10",X"20",X"00",X"FD",X"04",X"68",X"18",
		X"82",X"E7",X"20",X"6F",X"E7",X"50",X"03",X"20",
		X"82",X"E7",X"20",X"59",X"E7",X"56",X"50",X"4C",
		X"36",X"E7",X"FF",X"FF",X"C1",X"FF",X"7F",X"D1",
		X"CC",X"C7",X"CF",X"CE",X"C5",X"9A",X"98",X"8B",
		X"96",X"95",X"93",X"BF",X"B2",X"32",X"2D",X"2B",
		X"BC",X"B0",X"AC",X"BE",X"35",X"8E",X"61",X"FF",
		X"FF",X"FF",X"DD",X"FB",X"20",X"C9",X"EF",X"15",
		X"4F",X"10",X"05",X"20",X"C9",X"EF",X"35",X"4F",
		X"95",X"50",X"10",X"CB",X"4C",X"C9",X"EF",X"40",
		X"60",X"8D",X"60",X"8B",X"00",X"7E",X"8C",X"33",
		X"00",X"00",X"60",X"03",X"BF",X"12",X"00",X"40",
		X"89",X"C9",X"47",X"9D",X"17",X"68",X"9D",X"0A",
		X"00",X"40",X"60",X"8D",X"60",X"8B",X"00",X"7E",
		X"8C",X"3C",X"00",X"00",X"60",X"03",X"BF",X"1B",
		X"4B",X"67",X"B4",X"A1",X"07",X"8C",X"07",X"AE",
		X"A9",X"AC",X"A8",X"67",X"8C",X"07",X"B4",X"AF",
		X"AC",X"B0",X"67",X"9D",X"B2",X"AF",X"AC",X"AF",
		X"A3",X"67",X"8C",X"07",X"A5",X"AB",X"AF",X"B0",
		X"F4",X"AE",X"A9",X"B2",X"B0",X"7F",X"0E",X"27",
		X"B4",X"AE",X"A9",X"B2",X"B0",X"7F",X"0E",X"28",
		X"B4",X"AE",X"A9",X"B2",X"B0",X"64",X"07",X"A6",
		X"A9",X"67",X"AF",X"B4",X"AF",X"A7",X"78",X"B4",
		X"A5",X"AC",X"78",X"7F",X"02",X"AD",X"A5",X"B2",
		X"67",X"A2",X"B5",X"B3",X"AF",X"A7",X"EE",X"B2",
		X"B5",X"B4",X"A5",X"B2",X"7E",X"8C",X"39",X"B4",
		X"B8",X"A5",X"AE",X"67",X"B0",X"A5",X"B4",X"B3",
		X"27",X"AF",X"B4",X"07",X"9D",X"19",X"B2",X"AF",
		X"A6",X"7F",X"05",X"37",X"B4",X"B5",X"B0",X"AE",
		X"A9",X"7F",X"05",X"28",X"B4",X"B5",X"B0",X"AE",
		X"A9",X"7F",X"05",X"2A",X"B4",X"B5",X"B0",X"AE",
		X"A9",X"E4",X"AE",X"A5",X"ED",X"00",X"00",X"00",
		X"FF",X"FF",X"47",X"00",X"FD",X"04",X"68",X"18",
		X"A2",X"A1",X"B4",X"7F",X"0D",X"30",X"AD",X"A9",
		X"A4",X"7F",X"0D",X"23",X"AD",X"A9",X"A4",X"67",
		X"AC",X"AC",X"A1",X"A3",X"00",X"40",X"80",X"C0",
		X"C1",X"80",X"00",X"47",X"8C",X"68",X"8C",X"DB",
		X"67",X"9B",X"68",X"9B",X"50",X"8C",X"63",X"8C",
		X"7F",X"01",X"51",X"07",X"88",X"29",X"84",X"80",
		X"C4",X"80",X"57",X"71",X"07",X"88",X"14",X"ED",
		X"A5",X"AD",X"AF",X"AC",X"ED",X"A5",X"AD",X"A9",
		X"A8",X"F2",X"AF",X"AC",X"AF",X"A3",X"71",X"08",
		X"88",X"AE",X"A5",X"AC",X"68",X"83",X"08",X"68",
		X"9D",X"08",X"71",X"07",X"88",X"60",X"76",X"B4",
		X"AF",X"AE",X"76",X"8D",X"76",X"8B",X"51",X"07",
		X"88",X"19",X"B8",X"A4",X"AE",X"B2",X"F2",X"B3",
		X"B5",X"F3",X"A2",X"A1",X"EE",X"A7",X"B3",X"E4",
		X"AE",X"B2",X"EB",X"A5",X"A5",X"B0",X"51",X"07",
		X"88",X"39",X"81",X"C1",X"4F",X"7F",X"0F",X"2F",
		X"00",X"51",X"06",X"88",X"29",X"C2",X"0C",X"82",
		X"57",X"8C",X"6A",X"8C",X"42",X"AE",X"A5",X"A8",
		X"B4",X"60",X"AE",X"A5",X"A8",X"B4",X"4F",X"7E",
		X"1E",X"35",X"8C",X"27",X"51",X"07",X"88",X"09",
		X"8B",X"FE",X"E4",X"AF",X"AD",X"F2",X"AF",X"E4",
		X"AE",X"A1",X"DC",X"DE",X"9C",X"DD",X"9C",X"DE",
		X"DD",X"9E",X"C3",X"DD",X"CF",X"CA",X"CD",X"CB",
		X"00",X"47",X"9D",X"AD",X"A5",X"AD",X"AF",X"AC",
		X"76",X"9D",X"AD",X"A5",X"AD",X"A9",X"A8",X"E6",
		X"A6",X"AF",X"60",X"8C",X"20",X"AF",X"B4",X"B5",
		X"A1",X"F2",X"AC",X"A3",X"F2",X"A3",X"B3",X"60",
		X"8C",X"20",X"AC",X"A5",X"A4",X"EE",X"B5",X"B2",
		X"60",X"AE",X"B5",X"B2",X"F4",X"B3",X"A9",X"AC",
		X"60",X"8C",X"20",X"B4",X"B3",X"A9",X"AC",X"7A",
		X"7E",X"9A",X"22",X"20",X"00",X"60",X"03",X"BF",
		X"60",X"03",X"BF",X"00",X"FD",X"04",X"68",X"18",
		X"1F",X"EE",X"00",X"00",X"20",X"B1",X"E7",X"E8",
		X"E8",X"B5",X"4F",X"85",X"DA",X"B5",X"87",X"85",
		X"DB",X"B4",X"4E",X"98",X"D5",X"86",X"B0",X"09",
		X"B1",X"DA",X"20",X"C9",X"E3",X"C8",X"4C",X"0F",
		X"EE",X"A9",X"FF",X"85",X"D5",X"60",X"E8",X"A9",
		X"00",X"95",X"88",X"95",X"A8",X"B5",X"87",X"38",
		X"F5",X"4F",X"95",X"50",X"4C",X"23",X"E8",X"FF",
		X"20",X"15",X"E7",X"A5",X"CF",X"D0",X"28",X"A5",
		X"CE",X"60",X"20",X"34",X"EE",X"A4",X"C8",X"C9",
		X"30",X"B0",X"21",X"C0",X"28",X"B0",X"1D",X"60",
		X"EA",X"EA",X"20",X"34",X"EE",X"60",X"EA",X"8A",
		X"A2",X"01",X"B4",X"CE",X"94",X"4C",X"B4",X"48",
		X"94",X"CA",X"CA",X"F0",X"F5",X"AA",X"60",X"A0",
		X"77",X"4C",X"E0",X"E3",X"A0",X"7B",X"D0",X"F9",
		X"20",X"54",X"E2",X"A5",X"DA",X"D0",X"07",X"A5",
		X"DB",X"D0",X"03",X"4C",X"7E",X"E7",X"06",X"CE",
		X"26",X"CF",X"26",X"46",X"26",X"47",X"A5",X"46",
		X"C5",X"DA",X"A5",X"47",X"E5",X"DB",X"90",X"0A",
		X"85",X"47",X"A5",X"46",X"E5",X"DA",X"85",X"46",
		X"E6",X"CE",X"88",X"D0",X"E1",X"60",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"20",X"15",X"E7",X"6C",
		X"CE",X"00",X"A5",X"4C",X"D0",X"02",X"C6",X"4D",
		X"C6",X"4C",X"A5",X"48",X"D0",X"02",X"C6",X"49",
		X"C6",X"48",X"A0",X"00",X"B1",X"4C",X"91",X"48",
		X"A5",X"CA",X"C5",X"4C",X"A5",X"CB",X"E5",X"4D",
		X"90",X"E0",X"4C",X"53",X"EE",X"C9",X"28",X"B0",
		X"9B",X"A8",X"A5",X"C8",X"60",X"EA",X"EA",X"98",
		X"AA",X"A0",X"6E",X"20",X"C4",X"E3",X"8A",X"A8",
		X"20",X"C4",X"E3",X"A0",X"72",X"4C",X"C4",X"E3",
		X"20",X"15",X"E7",X"06",X"CE",X"26",X"CF",X"30",
		X"FA",X"B0",X"DC",X"D0",X"04",X"C5",X"CE",X"B0",
		X"D6",X"60",X"20",X"00",X"FD",X"04",X"68",X"18",
		X"15",X"E7",X"B1",X"CE",X"94",X"A7",X"4C",X"08",
		X"E7",X"EF",X"00",X"00",X"20",X"34",X"EE",X"A5",
		X"CE",X"48",X"20",X"15",X"E7",X"68",X"91",X"CE",
		X"60",X"FF",X"FF",X"FF",X"20",X"6C",X"EE",X"A5",
		X"CE",X"85",X"46",X"A5",X"CF",X"85",X"47",X"4C",
		X"44",X"E2",X"20",X"E4",X"EE",X"4C",X"34",X"E1",
		X"20",X"E4",X"EE",X"B4",X"88",X"B5",X"50",X"69",
		X"FE",X"B0",X"01",X"88",X"85",X"DA",X"84",X"DB",
		X"18",X"65",X"CE",X"95",X"50",X"98",X"65",X"CF",
		X"95",X"88",X"A0",X"00",X"B5",X"50",X"D1",X"DA",
		X"C8",X"B5",X"88",X"F1",X"DA",X"B0",X"80",X"4C",
		X"23",X"E8",X"20",X"15",X"E7",X"A5",X"4E",X"20",
		X"08",X"E7",X"A5",X"4F",X"D0",X"04",X"C5",X"4E",
		X"69",X"00",X"29",X"7F",X"85",X"4F",X"95",X"A8",
		X"A0",X"11",X"A5",X"4F",X"0A",X"18",X"69",X"40",
		X"0A",X"26",X"4E",X"26",X"4F",X"88",X"D0",X"F2",
		X"A5",X"CE",X"20",X"08",X"E7",X"A5",X"CF",X"95",
		X"A8",X"4C",X"7A",X"E2",X"20",X"15",X"E7",X"A4",
		X"CE",X"C4",X"4C",X"A5",X"CF",X"E5",X"4D",X"90",
		X"1F",X"84",X"48",X"A5",X"CF",X"85",X"49",X"4C",
		X"B6",X"EE",X"20",X"15",X"E7",X"A4",X"CE",X"C4",
		X"CA",X"A5",X"CF",X"E5",X"CB",X"B0",X"09",X"84",
		X"4A",X"A5",X"CF",X"85",X"4B",X"4C",X"B7",X"E5",
		X"4C",X"CB",X"EE",X"EA",X"EA",X"EA",X"EA",X"20",
		X"C9",X"EF",X"20",X"71",X"E1",X"4C",X"BF",X"EF",
		X"20",X"03",X"EE",X"A9",X"FF",X"85",X"C8",X"A9",
		X"74",X"8D",X"00",X"02",X"60",X"20",X"36",X"E7",
		X"E8",X"20",X"36",X"E7",X"B5",X"50",X"60",X"A9",
		X"00",X"85",X"4A",X"85",X"4C",X"A9",X"08",X"85",
		X"4B",X"A9",X"10",X"85",X"4D",X"4C",X"AD",X"E5",
		X"D5",X"88",X"D0",X"01",X"18",X"4C",X"02",X"E1",
		X"20",X"B7",X"E5",X"00",X"FD",X"04",X"68",X"18",
		X"4C",X"36",X"E8",X"20",X"B7",X"E5",X"4C",X"5B",
		X"E8",X"E0",X"80",X"D0",X"01",X"88",X"4C",X"0C",
		X"E0",X"FF",X"00",X"00",X"D8",X"58",X"A0",X"7F",
		X"8C",X"12",X"D0",X"A9",X"A7",X"8D",X"11",X"D0",
		X"8D",X"13",X"D0",X"C9",X"DF",X"F0",X"13",X"C9",
		X"9B",X"F0",X"03",X"C8",X"10",X"0F",X"A9",X"DC",
		X"20",X"EF",X"FF",X"A9",X"8D",X"20",X"EF",X"FF",
		X"A0",X"01",X"88",X"30",X"F6",X"AD",X"11",X"D0",
		X"10",X"FB",X"AD",X"10",X"D0",X"99",X"00",X"02",
		X"20",X"EF",X"FF",X"C9",X"8D",X"D0",X"D4",X"A0",
		X"FF",X"A9",X"00",X"AA",X"0A",X"85",X"3B",X"C8",
		X"B9",X"00",X"02",X"C9",X"8D",X"F0",X"D4",X"C9",
		X"AE",X"90",X"F4",X"F0",X"F0",X"C9",X"BA",X"F0",
		X"EB",X"C9",X"D2",X"F0",X"3B",X"86",X"38",X"86",
		X"39",X"84",X"3A",X"B9",X"00",X"02",X"49",X"B0",
		X"C9",X"0A",X"90",X"06",X"69",X"88",X"C9",X"FA",
		X"90",X"11",X"0A",X"0A",X"0A",X"0A",X"A2",X"04",
		X"0A",X"26",X"38",X"26",X"39",X"CA",X"D0",X"F8",
		X"C8",X"D0",X"E0",X"C4",X"3A",X"F0",X"97",X"24",
		X"3B",X"50",X"10",X"A5",X"38",X"81",X"36",X"E6",
		X"36",X"D0",X"B5",X"E6",X"37",X"4C",X"44",X"FF",
		X"6C",X"34",X"00",X"30",X"2B",X"A2",X"02",X"B5",
		X"37",X"95",X"35",X"95",X"33",X"CA",X"D0",X"F7",
		X"D0",X"14",X"A9",X"8D",X"20",X"EF",X"FF",X"A5",
		X"35",X"20",X"DC",X"FF",X"A5",X"34",X"20",X"DC",
		X"FF",X"A9",X"BA",X"20",X"EF",X"FF",X"A9",X"A0",
		X"20",X"EF",X"FF",X"A1",X"34",X"20",X"DC",X"FF",
		X"86",X"3B",X"A5",X"34",X"C5",X"38",X"A5",X"35",
		X"E5",X"39",X"B0",X"C1",X"E6",X"34",X"D0",X"02",
		X"E6",X"35",X"A5",X"34",X"29",X"07",X"10",X"C8",
		X"48",X"4A",X"4A",X"4A",X"4A",X"20",X"E5",X"FF",
		X"68",X"29",X"0F",X"00",X"FD",X"04",X"68",X"18",
		X"09",X"B0",X"C9",X"BA",X"90",X"02",X"69",X"06",
		X"8D",X"12",X"D0",X"2C",X"12",X"D0",X"D0",X"FB",
		X"60",X"00",X"00",X"00",X"00",X"00",X"FF",X"DB",
		X"5E",X"00",X"00",X"41",X"70",X"70",X"6C",X"65",
		X"31",X"00",X"00",X"8F",X"18",X"A2",X"FB",X"EE",
		X"19",X"02",X"00",X"12",X"1A",X"21",X"E6",X"38",
		X"35",X"53",X"0B",X"21",X"0E",X"F3",X"17",X"90",
		X"05",X"11",X"00",X"24",X"CF",X"18",X"02",X"18",
		X"E8",X"27",X"09",X"3E",X"08",X"90",X"0D",X"E6",
		X"09",X"51",X"0C",X"C5",X"10",X"7F",X"0C",X"93",
		X"0A",X"93",X"09",X"6B",X"09",X"16",X"0A",X"16",
		X"09",X"76",X"09",X"C0",X"09",X"29",X"0A",X"25",
		X"09",X"39",X"0A",X"71",X"18",X"FF",X"31",X"FF",
		X"2F",X"6D",X"0F",X"EE",X"13",X"68",X"18",X"78",
		X"0B",X"51",X"09",X"9B",X"07",X"5D",X"07",X"3F",
		X"0C",X"41",X"07",X"B1",X"1C",X"44",X"1D",X"D0",
		X"1C",X"38",X"00",X"B8",X"13",X"D9",X"13",X"CA",
		X"1F",X"EB",X"20",X"62",X"1A",X"46",X"20",X"40",
		X"21",X"47",X"21",X"90",X"21",X"FE",X"21",X"4A",
		X"18",X"B8",X"17",X"A1",X"14",X"E9",X"17",X"C7",
		X"17",X"28",X"17",X"3C",X"17",X"68",X"17",X"73",
		X"17",X"79",X"E1",X"18",X"79",X"97",X"18",X"7B",
		X"A2",X"1A",X"7B",X"89",X"1B",X"7F",X"D3",X"1F",
		X"50",X"2D",X"10",X"46",X"2A",X"10",X"7D",X"0C",
		X"20",X"5A",X"39",X"0F",X"64",X"5A",X"10",X"45",
		X"4E",X"C4",X"46",X"4F",X"D2",X"4E",X"45",X"58",
		X"D4",X"44",X"41",X"54",X"C1",X"49",X"4E",X"50",
		X"55",X"D4",X"44",X"49",X"CD",X"52",X"45",X"41",
		X"C4",X"4C",X"45",X"D4",X"47",X"4F",X"54",X"CF",
		X"52",X"55",X"CE",X"49",X"C6",X"52",X"45",X"53",
		X"54",X"4F",X"52",X"C5",X"47",X"4F",X"53",X"55",
		X"C2",X"52",X"45",X"00",X"FD",X"04",X"68",X"18",
		X"54",X"55",X"52",X"CE",X"52",X"45",X"CD",X"53",
		X"54",X"4F",X"D0",X"4F",X"CE",X"57",X"41",X"49",
		X"D4",X"4C",X"4F",X"41",X"C4",X"53",X"41",X"56",
		X"C5",X"56",X"45",X"52",X"49",X"46",X"D9",X"44",
		X"45",X"C6",X"50",X"4F",X"4B",X"C5",X"50",X"52",
		X"49",X"4E",X"D4",X"43",X"4F",X"4E",X"03",X"00",
		X"00",X"D4",X"4C",X"49",X"53",X"D4",X"43",X"4C",
		X"D2",X"47",X"45",X"D4",X"4E",X"45",X"D7",X"54",
		X"41",X"42",X"A8",X"54",X"CF",X"46",X"CE",X"53",
		X"50",X"43",X"A8",X"54",X"48",X"45",X"CE",X"4E",
		X"4F",X"D4",X"53",X"54",X"45",X"D0",X"AB",X"AD",
		X"AA",X"AF",X"DE",X"41",X"4E",X"C4",X"4F",X"D2",
		X"BE",X"BD",X"BC",X"53",X"47",X"CE",X"49",X"4E",
		X"D4",X"41",X"42",X"D3",X"55",X"53",X"D2",X"46",
		X"52",X"C5",X"50",X"4F",X"D3",X"53",X"51",X"D2",
		X"52",X"4E",X"C4",X"4C",X"4F",X"C7",X"45",X"58",
		X"D0",X"43",X"4F",X"D3",X"53",X"49",X"CE",X"54",
		X"41",X"CE",X"41",X"54",X"CE",X"50",X"45",X"45",
		X"CB",X"4C",X"45",X"CE",X"53",X"54",X"52",X"A4",
		X"56",X"41",X"CC",X"41",X"53",X"C3",X"43",X"48",
		X"52",X"A4",X"4C",X"45",X"46",X"54",X"A4",X"52",
		X"49",X"47",X"48",X"54",X"A4",X"4D",X"49",X"44",
		X"A4",X"47",X"CF",X"00",X"4E",X"45",X"58",X"54",
		X"20",X"57",X"49",X"54",X"48",X"4F",X"55",X"54",
		X"20",X"46",X"4F",X"D2",X"53",X"59",X"4E",X"54",
		X"41",X"D8",X"52",X"45",X"54",X"55",X"52",X"4E",
		X"20",X"57",X"49",X"54",X"48",X"4F",X"55",X"54",
		X"20",X"47",X"4F",X"53",X"55",X"C2",X"4F",X"55",
		X"54",X"20",X"4F",X"46",X"20",X"44",X"41",X"54",
		X"C1",X"49",X"4C",X"4C",X"45",X"47",X"41",X"4C",
		X"20",X"51",X"55",X"41",X"4E",X"54",X"49",X"54",
		X"D9",X"4F",X"56",X"00",X"FD",X"04",X"68",X"18",
		X"45",X"52",X"46",X"4C",X"4F",X"D7",X"4F",X"55",
		X"54",X"20",X"4F",X"46",X"20",X"4D",X"45",X"4D",
		X"4F",X"52",X"D9",X"55",X"4E",X"44",X"45",X"46",
		X"27",X"44",X"20",X"53",X"54",X"41",X"54",X"45",
		X"4D",X"45",X"4E",X"D4",X"42",X"41",X"44",X"20",
		X"53",X"55",X"42",X"53",X"43",X"52",X"49",X"50",
		X"D4",X"52",X"45",X"44",X"49",X"4D",X"04",X"00",
		X"00",X"27",X"44",X"20",X"41",X"52",X"52",X"41",
		X"D9",X"44",X"49",X"56",X"49",X"53",X"49",X"4F",
		X"4E",X"20",X"42",X"59",X"20",X"5A",X"45",X"52",
		X"CF",X"49",X"4C",X"4C",X"45",X"47",X"41",X"4C",
		X"20",X"44",X"49",X"52",X"45",X"43",X"D4",X"54",
		X"59",X"50",X"45",X"20",X"4D",X"49",X"53",X"4D",
		X"41",X"54",X"43",X"C8",X"53",X"54",X"52",X"49",
		X"4E",X"47",X"20",X"54",X"4F",X"4F",X"20",X"4C",
		X"4F",X"4E",X"C7",X"46",X"4F",X"52",X"4D",X"55",
		X"4C",X"41",X"20",X"54",X"4F",X"4F",X"20",X"43",
		X"4F",X"4D",X"50",X"4C",X"45",X"D8",X"43",X"41",
		X"4E",X"27",X"54",X"20",X"43",X"4F",X"4E",X"54",
		X"49",X"4E",X"55",X"C5",X"55",X"4E",X"44",X"45",
		X"46",X"27",X"44",X"20",X"46",X"55",X"4E",X"43",
		X"54",X"49",X"4F",X"CE",X"20",X"00",X"2E",X"38",
		X"4C",X"CC",X"0F",X"A0",X"1B",X"18",X"88",X"69",
		X"06",X"90",X"FB",X"60",X"20",X"45",X"52",X"52",
		X"4F",X"52",X"00",X"20",X"49",X"4E",X"20",X"00",
		X"0D",X"0A",X"52",X"45",X"41",X"44",X"59",X"2E",
		X"0D",X"0A",X"00",X"0D",X"0A",X"42",X"52",X"45",
		X"41",X"4B",X"00",X"BA",X"E8",X"E8",X"E8",X"E8",
		X"B5",X"01",X"C9",X"81",X"D0",X"1D",X"A5",X"7C",
		X"D0",X"08",X"B5",X"02",X"85",X"7B",X"B5",X"03",
		X"85",X"7C",X"D5",X"03",X"D0",X"06",X"A5",X"7B",
		X"D5",X"02",X"F0",X"00",X"FD",X"04",X"68",X"18",
		X"07",X"8A",X"18",X"69",X"12",X"AA",X"D0",X"DD",
		X"60",X"20",X"1B",X"05",X"85",X"63",X"84",X"64",
		X"38",X"A5",X"8D",X"E5",X"92",X"85",X"54",X"A8",
		X"A5",X"8E",X"E5",X"93",X"AA",X"E8",X"98",X"F0",
		X"23",X"A5",X"8D",X"38",X"E5",X"54",X"85",X"8D",
		X"B0",X"03",X"C6",X"8E",X"38",X"A5",X"8B",X"E5",
		X"54",X"85",X"8B",X"B0",X"08",X"C6",X"8C",X"90",
		X"04",X"B1",X"8D",X"91",X"8B",X"88",X"05",X"00",
		X"00",X"D0",X"F9",X"B1",X"8D",X"91",X"8B",X"C6",
		X"8E",X"C6",X"8C",X"CA",X"D0",X"F2",X"60",X"0A",
		X"69",X"B2",X"B0",X"35",X"85",X"54",X"BA",X"E4",
		X"54",X"90",X"2E",X"60",X"C4",X"66",X"90",X"28",
		X"D0",X"04",X"C5",X"65",X"90",X"22",X"48",X"A2",
		X"09",X"98",X"48",X"B5",X"8A",X"CA",X"10",X"FA",
		X"20",X"62",X"15",X"A2",X"F7",X"68",X"95",X"94",
		X"E8",X"30",X"FA",X"68",X"A8",X"68",X"C4",X"66",
		X"90",X"06",X"D0",X"05",X"C5",X"65",X"B0",X"01",
		X"60",X"A2",X"4D",X"46",X"45",X"20",X"AC",X"0B",
		X"20",X"0F",X"0C",X"BD",X"83",X"03",X"48",X"29",
		X"7F",X"20",X"11",X"0C",X"E8",X"68",X"10",X"F3",
		X"20",X"7A",X"07",X"A9",X"83",X"A0",X"04",X"20",
		X"EF",X"0B",X"A4",X"6C",X"C8",X"F0",X"03",X"20",
		X"3A",X"1E",X"46",X"45",X"A9",X"8F",X"A0",X"04",
		X"20",X"EF",X"0B",X"20",X"57",X"06",X"86",X"A6",
		X"84",X"A7",X"20",X"6B",X"22",X"AA",X"F0",X"F3",
		X"A2",X"FF",X"86",X"6C",X"90",X"06",X"20",X"7E",
		X"06",X"4C",X"DE",X"08",X"20",X"5A",X"0A",X"20",
		X"7E",X"06",X"84",X"3D",X"20",X"13",X"07",X"90",
		X"44",X"A0",X"01",X"B1",X"92",X"85",X"55",X"A5",
		X"5F",X"85",X"54",X"A5",X"93",X"85",X"57",X"A5",
		X"92",X"88",X"F1",X"92",X"18",X"65",X"5F",X"85",
		X"5F",X"85",X"56",X"00",X"FD",X"04",X"68",X"18",
		X"A5",X"60",X"69",X"FF",X"85",X"60",X"E5",X"93",
		X"AA",X"38",X"A5",X"92",X"E5",X"5F",X"A8",X"B0",
		X"03",X"E8",X"C6",X"57",X"18",X"65",X"54",X"90",
		X"03",X"C6",X"55",X"18",X"B1",X"54",X"91",X"56",
		X"C8",X"D0",X"F9",X"E6",X"55",X"E6",X"57",X"CA",
		X"D0",X"F2",X"20",X"59",X"07",X"20",X"2A",X"06",
		X"AD",X"05",X"24",X"F0",X"8B",X"18",X"A5",X"5F",
		X"85",X"8D",X"65",X"3D",X"85",X"8B",X"A4",X"60",
		X"84",X"8E",X"90",X"01",X"C8",X"84",X"06",X"00",
		X"00",X"8C",X"20",X"CB",X"04",X"A5",X"46",X"A4",
		X"47",X"8D",X"03",X"24",X"8C",X"04",X"24",X"A5",
		X"63",X"A4",X"64",X"85",X"5F",X"84",X"60",X"A4",
		X"3D",X"88",X"B9",X"01",X"24",X"91",X"92",X"88",
		X"10",X"F8",X"20",X"59",X"07",X"20",X"2A",X"06",
		X"4C",X"7A",X"05",X"A5",X"5D",X"A4",X"5E",X"85",
		X"54",X"84",X"55",X"18",X"A0",X"01",X"B1",X"54",
		X"F0",X"1D",X"A0",X"04",X"C8",X"B1",X"54",X"D0",
		X"FB",X"C8",X"98",X"65",X"54",X"AA",X"A0",X"00",
		X"91",X"54",X"A5",X"55",X"69",X"00",X"C8",X"91",
		X"54",X"86",X"54",X"85",X"55",X"90",X"DD",X"60",
		X"A2",X"00",X"20",X"6E",X"06",X"C9",X"0D",X"F0",
		X"0B",X"20",X"00",X"2F",X"F0",X"F4",X"9D",X"05",
		X"24",X"E8",X"D0",X"EE",X"4C",X"A3",X"0B",X"20",
		X"00",X"2C",X"C9",X"0F",X"D0",X"08",X"48",X"A5",
		X"45",X"49",X"FF",X"85",X"45",X"68",X"60",X"A6",
		X"A6",X"A0",X"04",X"84",X"41",X"BD",X"00",X"24",
		X"10",X"07",X"C9",X"FF",X"F0",X"3E",X"E8",X"D0",
		X"F4",X"C9",X"20",X"F0",X"37",X"85",X"3C",X"C9",
		X"22",X"F0",X"56",X"24",X"41",X"70",X"2D",X"C9",
		X"3F",X"D0",X"04",X"A9",X"97",X"D0",X"25",X"C9",
		X"30",X"90",X"04",X"C9",X"3C",X"90",X"1D",X"84",
		X"A4",X"A0",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"84",X"3D",X"88",X"86",X"A6",X"CA",X"C8",X"E8",
		X"BD",X"00",X"24",X"38",X"F9",X"9E",X"02",X"F0",
		X"F5",X"C9",X"80",X"D0",X"30",X"05",X"3D",X"A4",
		X"A4",X"E8",X"C8",X"99",X"00",X"24",X"B9",X"00",
		X"24",X"F0",X"36",X"38",X"E9",X"3A",X"F0",X"04",
		X"C9",X"49",X"D0",X"02",X"85",X"41",X"38",X"E9",
		X"54",X"D0",X"9F",X"85",X"3C",X"BD",X"00",X"24",
		X"F0",X"DF",X"C5",X"3C",X"F0",X"DB",X"C8",X"99",
		X"00",X"24",X"E8",X"D0",X"F0",X"A6",X"A6",X"E6",
		X"3D",X"C8",X"B9",X"9D",X"02",X"10",X"07",X"00",
		X"00",X"FA",X"B9",X"9E",X"02",X"D0",X"B4",X"BD",
		X"00",X"24",X"10",X"BE",X"99",X"02",X"24",X"A9",
		X"04",X"85",X"A6",X"60",X"A5",X"5D",X"A6",X"5E",
		X"A0",X"01",X"85",X"92",X"86",X"93",X"B1",X"92",
		X"F0",X"1F",X"C8",X"C8",X"A5",X"47",X"D1",X"92",
		X"90",X"18",X"F0",X"03",X"88",X"D0",X"09",X"A5",
		X"46",X"88",X"D1",X"92",X"90",X"0C",X"F0",X"0A",
		X"88",X"B1",X"92",X"AA",X"88",X"B1",X"92",X"B0",
		X"D7",X"18",X"60",X"D0",X"FD",X"A9",X"00",X"A8",
		X"91",X"5D",X"C8",X"91",X"5D",X"A5",X"5D",X"18",
		X"69",X"02",X"85",X"5F",X"A5",X"5E",X"69",X"00",
		X"85",X"60",X"20",X"8E",X"07",X"A9",X"00",X"D0",
		X"2D",X"A5",X"69",X"A4",X"6A",X"85",X"65",X"84",
		X"66",X"20",X"00",X"2E",X"A5",X"5F",X"A4",X"60",
		X"85",X"61",X"84",X"62",X"85",X"63",X"84",X"64",
		X"20",X"17",X"09",X"A2",X"4B",X"86",X"48",X"68",
		X"A8",X"68",X"A2",X"FF",X"9A",X"48",X"98",X"48",
		X"A9",X"00",X"85",X"70",X"85",X"42",X"60",X"18",
		X"A5",X"5D",X"69",X"FF",X"85",X"A6",X"A5",X"5E",
		X"69",X"FF",X"85",X"A7",X"60",X"90",X"06",X"F0",
		X"04",X"C9",X"A5",X"D0",X"E9",X"20",X"5A",X"0A",
		X"20",X"13",X"07",X"00",X"FD",X"04",X"68",X"18",
		X"20",X"71",X"22",X"F0",X"0C",X"C9",X"A5",X"D0",
		X"8E",X"20",X"6B",X"22",X"20",X"5A",X"0A",X"D0",
		X"86",X"68",X"68",X"A5",X"46",X"05",X"47",X"D0",
		X"06",X"A9",X"FF",X"85",X"46",X"85",X"47",X"A0",
		X"01",X"84",X"41",X"B1",X"92",X"F0",X"43",X"20",
		X"00",X"2D",X"20",X"AC",X"0B",X"C8",X"B1",X"92",
		X"AA",X"C8",X"B1",X"92",X"C5",X"47",X"D0",X"04",
		X"E4",X"46",X"F0",X"02",X"B0",X"2C",X"84",X"7B",
		X"20",X"45",X"1E",X"A9",X"20",X"A4",X"7B",X"29",
		X"7F",X"20",X"11",X"0C",X"C9",X"22",X"D0",X"06",
		X"A5",X"41",X"49",X"FF",X"85",X"41",X"08",X"00",
		X"00",X"C8",X"F0",X"11",X"B1",X"92",X"D0",X"10",
		X"A8",X"B1",X"92",X"AA",X"C8",X"B1",X"92",X"86",
		X"92",X"85",X"93",X"D0",X"B5",X"4C",X"71",X"05",
		X"10",X"DA",X"C9",X"FF",X"F0",X"D6",X"24",X"41",
		X"30",X"D2",X"38",X"E9",X"7F",X"AA",X"84",X"7B",
		X"A0",X"FF",X"CA",X"F0",X"08",X"C8",X"B9",X"9E",
		X"02",X"10",X"FA",X"30",X"F5",X"C8",X"B9",X"9E",
		X"02",X"30",X"B5",X"20",X"11",X"0C",X"D0",X"F5",
		X"A9",X"80",X"85",X"42",X"20",X"94",X"0A",X"20",
		X"A2",X"04",X"D0",X"05",X"8A",X"69",X"0F",X"AA",
		X"9A",X"68",X"68",X"A9",X"09",X"20",X"0E",X"05",
		X"20",X"F5",X"09",X"18",X"98",X"65",X"A6",X"48",
		X"A5",X"A7",X"69",X"00",X"48",X"A5",X"6C",X"48",
		X"A5",X"6B",X"48",X"A9",X"9E",X"20",X"65",X"0F",
		X"20",X"F9",X"0D",X"20",X"F6",X"0D",X"A5",X"99",
		X"09",X"7F",X"25",X"95",X"85",X"95",X"A9",X"88",
		X"A0",X"08",X"85",X"54",X"84",X"55",X"4C",X"AF",
		X"0E",X"A9",X"34",X"A0",X"1A",X"20",X"1A",X"1C",
		X"20",X"71",X"22",X"C9",X"A3",X"D0",X"06",X"20",
		X"6B",X"22",X"20",X"F6",X"0D",X"20",X"A3",X"1C",
		X"20",X"A4",X"0E",X"00",X"FD",X"04",X"68",X"18",
		X"A5",X"7C",X"48",X"A5",X"7B",X"48",X"A9",X"81",
		X"48",X"20",X"00",X"2D",X"A5",X"A6",X"A4",X"A7",
		X"C0",X"24",X"EA",X"F0",X"04",X"85",X"6F",X"84",
		X"70",X"A0",X"00",X"B1",X"A6",X"D0",X"40",X"A0",
		X"02",X"B1",X"A6",X"18",X"D0",X"03",X"4C",X"42",
		X"09",X"C8",X"B1",X"A6",X"85",X"6B",X"C8",X"B1",
		X"A6",X"85",X"6C",X"98",X"65",X"A6",X"85",X"A6",
		X"90",X"02",X"E6",X"A7",X"20",X"6B",X"22",X"20",
		X"E7",X"08",X"4C",X"AB",X"08",X"F0",X"3C",X"E9",
		X"80",X"90",X"11",X"C9",X"1D",X"B0",X"17",X"0A",
		X"A8",X"B9",X"19",X"02",X"48",X"B9",X"18",X"02",
		X"48",X"4C",X"6B",X"22",X"4C",X"94",X"09",X"00",
		X"00",X"0A",X"C9",X"3A",X"F0",X"D9",X"4C",X"6E",
		X"0F",X"C9",X"45",X"D0",X"F9",X"20",X"6B",X"22",
		X"A9",X"9E",X"20",X"65",X"0F",X"4C",X"94",X"09",
		X"38",X"A5",X"5D",X"E9",X"01",X"A4",X"5E",X"B0",
		X"01",X"88",X"85",X"73",X"84",X"74",X"60",X"B0",
		X"01",X"18",X"D0",X"40",X"A5",X"A6",X"A4",X"A7",
		X"A6",X"6C",X"E8",X"F0",X"0C",X"85",X"6F",X"84",
		X"70",X"A5",X"6B",X"A4",X"6C",X"85",X"6D",X"84",
		X"6E",X"68",X"68",X"A9",X"9A",X"A0",X"04",X"A2",
		X"00",X"86",X"45",X"90",X"03",X"4C",X"66",X"05",
		X"4C",X"71",X"05",X"D0",X"17",X"A2",X"D2",X"A4",
		X"70",X"D0",X"03",X"4C",X"4A",X"05",X"A5",X"6F",
		X"85",X"A6",X"84",X"A7",X"A5",X"6D",X"A4",X"6E",
		X"85",X"6B",X"84",X"6C",X"60",X"D0",X"03",X"4C",
		X"59",X"07",X"20",X"60",X"07",X"4C",X"8B",X"09",
		X"A9",X"03",X"20",X"0E",X"05",X"A5",X"A7",X"48",
		X"A5",X"A6",X"48",X"A5",X"6C",X"48",X"A5",X"6B",
		X"48",X"A9",X"8C",X"48",X"20",X"71",X"22",X"20",
		X"94",X"09",X"4C",X"AB",X"08",X"20",X"5A",X"0A",
		X"20",X"F8",X"09",X"00",X"FD",X"04",X"68",X"18",
		X"A5",X"6C",X"C5",X"47",X"B0",X"0B",X"98",X"38",
		X"65",X"A6",X"A6",X"A7",X"90",X"07",X"E8",X"B0",
		X"04",X"A5",X"5D",X"A6",X"5E",X"20",X"17",X"07",
		X"90",X"1E",X"A5",X"92",X"E9",X"01",X"85",X"A6",
		X"A5",X"93",X"E9",X"00",X"85",X"A7",X"60",X"D0",
		X"FD",X"A9",X"FF",X"85",X"7C",X"20",X"A2",X"04",
		X"9A",X"C9",X"8C",X"F0",X"0B",X"A2",X"16",X"2C",
		X"A2",X"5A",X"4C",X"4A",X"05",X"4C",X"6E",X"0F",
		X"68",X"68",X"85",X"6B",X"68",X"85",X"6C",X"68",
		X"85",X"A6",X"68",X"85",X"A7",X"20",X"F5",X"09",
		X"98",X"18",X"65",X"A6",X"85",X"A6",X"90",X"02",
		X"E6",X"A7",X"60",X"A2",X"3A",X"2C",X"A2",X"00",
		X"86",X"3B",X"A0",X"00",X"84",X"3C",X"0A",X"00",
		X"00",X"A5",X"3C",X"A6",X"3B",X"85",X"3B",X"86",
		X"3C",X"B1",X"A6",X"F0",X"E8",X"C5",X"3C",X"F0",
		X"E4",X"C8",X"C9",X"22",X"D0",X"F3",X"F0",X"E9",
		X"20",X"0A",X"0E",X"20",X"71",X"22",X"C9",X"88",
		X"F0",X"05",X"A9",X"A1",X"20",X"65",X"0F",X"A5",
		X"94",X"D0",X"05",X"20",X"F8",X"09",X"F0",X"BB",
		X"20",X"71",X"22",X"B0",X"03",X"4C",X"94",X"09",
		X"4C",X"E7",X"08",X"20",X"DA",X"17",X"48",X"C9",
		X"8C",X"F0",X"04",X"C9",X"88",X"D0",X"91",X"C6",
		X"98",X"D0",X"04",X"68",X"4C",X"E9",X"08",X"20",
		X"6B",X"22",X"20",X"5A",X"0A",X"C9",X"2C",X"F0",
		X"EE",X"68",X"60",X"A2",X"00",X"86",X"46",X"86",
		X"47",X"B0",X"F7",X"E9",X"2F",X"85",X"3B",X"A5",
		X"47",X"85",X"54",X"C9",X"19",X"B0",X"D4",X"A5",
		X"46",X"0A",X"26",X"54",X"0A",X"26",X"54",X"65",
		X"46",X"85",X"46",X"A5",X"54",X"65",X"47",X"85",
		X"47",X"06",X"46",X"26",X"47",X"A5",X"46",X"65",
		X"3B",X"85",X"46",X"90",X"02",X"E6",X"47",X"20",
		X"6B",X"22",X"4C",X"00",X"FD",X"04",X"68",X"18",
		X"60",X"0A",X"20",X"D0",X"10",X"85",X"7B",X"84",
		X"7C",X"A9",X"AC",X"20",X"65",X"0F",X"A5",X"40",
		X"48",X"A5",X"3F",X"48",X"20",X"0A",X"0E",X"68",
		X"2A",X"20",X"FC",X"0D",X"D0",X"18",X"68",X"10",
		X"12",X"20",X"93",X"1C",X"20",X"FD",X"11",X"A0",
		X"00",X"A5",X"97",X"91",X"7B",X"C8",X"A5",X"98",
		X"91",X"7B",X"60",X"4C",X"48",X"1C",X"68",X"A4",
		X"7C",X"C0",X"1F",X"D0",X"50",X"20",X"E2",X"16",
		X"C9",X"06",X"D0",X"41",X"A0",X"00",X"84",X"94",
		X"84",X"99",X"84",X"A4",X"20",X"10",X"0B",X"20",
		X"5A",X"1B",X"E6",X"A4",X"A4",X"A4",X"20",X"10",
		X"0B",X"20",X"84",X"1C",X"AA",X"F0",X"05",X"E8",
		X"8A",X"20",X"65",X"1B",X"A4",X"A4",X"C8",X"C0",
		X"06",X"D0",X"DF",X"20",X"5A",X"1B",X"0B",X"00",
		X"00",X"20",X"13",X"1D",X"A2",X"02",X"78",X"B5",
		X"96",X"9D",X"00",X"02",X"CA",X"10",X"F8",X"58",
		X"60",X"B1",X"54",X"20",X"7D",X"22",X"90",X"03",
		X"4C",X"82",X"12",X"E9",X"2F",X"4C",X"F6",X"1D",
		X"A0",X"02",X"B1",X"97",X"C5",X"66",X"90",X"17",
		X"D0",X"07",X"88",X"B1",X"97",X"C5",X"65",X"90",
		X"0E",X"A4",X"98",X"C4",X"60",X"90",X"08",X"D0",
		X"0D",X"A5",X"97",X"C5",X"5F",X"B0",X"07",X"A5",
		X"97",X"A4",X"98",X"4C",X"5B",X"0B",X"A0",X"00",
		X"B1",X"97",X"20",X"B1",X"14",X"A5",X"83",X"A4",
		X"84",X"85",X"A2",X"84",X"A3",X"20",X"B6",X"16",
		X"A9",X"94",X"A0",X"00",X"85",X"83",X"84",X"84",
		X"20",X"17",X"17",X"A0",X"00",X"B1",X"83",X"91",
		X"7B",X"C8",X"B1",X"83",X"91",X"7B",X"C8",X"B1",
		X"83",X"91",X"7B",X"60",X"20",X"F2",X"0B",X"20",
		X"71",X"22",X"F0",X"31",X"F0",X"3B",X"C9",X"9D",
		X"F0",X"49",X"C9",X"A0",X"18",X"F0",X"44",X"C9",
		X"2C",X"F0",X"2F",X"00",X"FD",X"04",X"68",X"18",
		X"C9",X"3B",X"F0",X"56",X"20",X"0A",X"0E",X"24",
		X"3F",X"30",X"DE",X"20",X"55",X"1E",X"20",X"C3",
		X"14",X"20",X"F2",X"0B",X"20",X"0C",X"0C",X"D0",
		X"D3",X"A9",X"00",X"9D",X"05",X"24",X"A2",X"04",
		X"A0",X"24",X"A9",X"0D",X"20",X"11",X"0C",X"A9",
		X"0A",X"20",X"11",X"0C",X"49",X"FF",X"60",X"A5",
		X"30",X"20",X"7A",X"04",X"98",X"38",X"E9",X"0A",
		X"B0",X"FC",X"49",X"FF",X"69",X"01",X"D0",X"15",
		X"08",X"20",X"D7",X"17",X"C9",X"29",X"D0",X"5B",
		X"28",X"90",X"0B",X"A5",X"30",X"20",X"7A",X"04",
		X"8A",X"E5",X"2B",X"90",X"05",X"AA",X"E8",X"CA",
		X"D0",X"06",X"20",X"6B",X"22",X"4C",X"7B",X"0B",
		X"20",X"0C",X"0C",X"D0",X"F2",X"20",X"C3",X"14",
		X"20",X"E2",X"16",X"AA",X"A0",X"00",X"E8",X"CA",
		X"F0",X"BC",X"B1",X"54",X"20",X"11",X"0C",X"00",
		X"00",X"0C",X"C8",X"C9",X"0D",X"D0",X"F3",X"20",
		X"B6",X"0B",X"4C",X"F9",X"0B",X"A9",X"20",X"2C",
		X"A9",X"3F",X"24",X"45",X"30",X"03",X"20",X"00",
		X"2B",X"29",X"FF",X"60",X"A5",X"43",X"F0",X"11",
		X"30",X"04",X"A0",X"FF",X"D0",X"04",X"A5",X"71",
		X"A4",X"72",X"85",X"6B",X"84",X"6C",X"4C",X"6E",
		X"0F",X"A9",X"7E",X"A0",X"0D",X"20",X"EF",X"0B",
		X"A5",X"6F",X"A4",X"70",X"85",X"A6",X"84",X"A7",
		X"60",X"20",X"E2",X"13",X"A2",X"06",X"A0",X"24",
		X"A9",X"00",X"8D",X"06",X"24",X"A9",X"40",X"20",
		X"89",X"0C",X"60",X"46",X"45",X"C9",X"22",X"D0",
		X"0B",X"20",X"23",X"0F",X"A9",X"3B",X"20",X"65",
		X"0F",X"20",X"F2",X"0B",X"20",X"E2",X"13",X"A9",
		X"2C",X"8D",X"04",X"24",X"20",X"77",X"0C",X"AD",
		X"05",X"24",X"D0",X"14",X"18",X"4C",X"38",X"09",
		X"20",X"0F",X"0C",X"20",X"0C",X"0C",X"4C",X"57",
		X"06",X"A6",X"73",X"00",X"FD",X"04",X"68",X"18",
		X"A4",X"74",X"A9",X"98",X"2C",X"A9",X"00",X"85",
		X"43",X"86",X"75",X"84",X"76",X"20",X"D0",X"10",
		X"85",X"7B",X"84",X"7C",X"A5",X"A6",X"A4",X"A7",
		X"85",X"7D",X"84",X"7E",X"A6",X"75",X"A4",X"76",
		X"86",X"A6",X"84",X"A7",X"20",X"71",X"22",X"D0",
		X"1C",X"24",X"43",X"50",X"0C",X"20",X"00",X"2C",
		X"8D",X"05",X"24",X"A2",X"04",X"A0",X"24",X"D0",
		X"08",X"30",X"71",X"20",X"0F",X"0C",X"20",X"77",
		X"0C",X"86",X"A6",X"84",X"A7",X"20",X"6B",X"22",
		X"24",X"3F",X"10",X"31",X"24",X"43",X"50",X"09",
		X"E8",X"86",X"A6",X"A9",X"00",X"85",X"3B",X"F0",
		X"0C",X"85",X"3B",X"C9",X"22",X"F0",X"07",X"A9",
		X"3A",X"85",X"3B",X"A9",X"2C",X"18",X"85",X"3C",
		X"A5",X"A6",X"A4",X"A7",X"69",X"00",X"90",X"01",
		X"C8",X"20",X"C9",X"14",X"20",X"1F",X"18",X"20",
		X"C9",X"0A",X"4C",X"07",X"0D",X"20",X"0D",X"00",
		X"00",X"6B",X"1D",X"A5",X"40",X"20",X"B1",X"0A",
		X"20",X"71",X"22",X"F0",X"07",X"C9",X"2C",X"F0",
		X"03",X"4C",X"1B",X"0C",X"A5",X"A6",X"A4",X"A7",
		X"85",X"75",X"84",X"76",X"A5",X"7D",X"A4",X"7E",
		X"85",X"A6",X"84",X"A7",X"20",X"71",X"22",X"F0",
		X"2C",X"20",X"63",X"0F",X"4C",X"8F",X"0C",X"20",
		X"F5",X"09",X"C8",X"AA",X"D0",X"12",X"A2",X"2A",
		X"C8",X"B1",X"A6",X"F0",X"69",X"C8",X"B1",X"A6",
		X"85",X"71",X"C8",X"B1",X"A6",X"C8",X"85",X"72",
		X"B1",X"A6",X"AA",X"20",X"EA",X"09",X"E0",X"83",
		X"D0",X"DD",X"4C",X"C7",X"0C",X"A5",X"75",X"A4",
		X"76",X"A6",X"43",X"10",X"03",X"4C",X"21",X"09",
		X"A0",X"00",X"B1",X"75",X"F0",X"07",X"A9",X"6D",
		X"A0",X"0D",X"4C",X"EF",X"0B",X"60",X"3F",X"45",
		X"58",X"54",X"52",X"41",X"20",X"49",X"47",X"4E",
		X"4F",X"52",X"45",X"00",X"FD",X"04",X"68",X"18",
		X"44",X"0D",X"0A",X"00",X"3F",X"52",X"45",X"44",
		X"4F",X"20",X"46",X"52",X"4F",X"4D",X"20",X"53",
		X"54",X"41",X"52",X"54",X"0D",X"0A",X"00",X"D0",
		X"04",X"A0",X"00",X"F0",X"03",X"20",X"D0",X"10",
		X"85",X"7B",X"84",X"7C",X"20",X"A2",X"04",X"F0",
		X"04",X"A2",X"00",X"F0",X"60",X"9A",X"8A",X"18",
		X"69",X"04",X"48",X"69",X"06",X"85",X"56",X"68",
		X"A0",X"00",X"20",X"1A",X"1C",X"BA",X"B5",X"09",
		X"85",X"99",X"A5",X"7B",X"A4",X"7C",X"20",X"DF",
		X"18",X"20",X"48",X"1C",X"A0",X"00",X"20",X"D5",
		X"1C",X"BA",X"38",X"F5",X"09",X"F0",X"13",X"B5",
		X"0F",X"85",X"6B",X"B5",X"10",X"85",X"6C",X"B5",
		X"12",X"85",X"A6",X"B5",X"11",X"85",X"A7",X"4C",
		X"AB",X"08",X"8A",X"69",X"11",X"AA",X"9A",X"20",
		X"71",X"22",X"C9",X"2C",X"D0",X"F1",X"20",X"6B",
		X"22",X"20",X"97",X"0D",X"20",X"0A",X"0E",X"18",
		X"24",X"38",X"24",X"3F",X"30",X"03",X"0E",X"00",
		X"00",X"B0",X"03",X"60",X"B0",X"FD",X"A2",X"A3",
		X"4C",X"4A",X"05",X"A6",X"A6",X"D0",X"02",X"C6",
		X"A7",X"C6",X"A6",X"A2",X"00",X"24",X"48",X"8A",
		X"48",X"A9",X"01",X"20",X"0E",X"05",X"20",X"EF",
		X"0E",X"A9",X"00",X"85",X"7F",X"20",X"71",X"22",
		X"38",X"E9",X"AB",X"90",X"17",X"C9",X"03",X"B0",
		X"13",X"C9",X"01",X"2A",X"49",X"01",X"45",X"7F",
		X"C5",X"7F",X"90",X"61",X"85",X"7F",X"20",X"6B",
		X"22",X"4C",X"27",X"0E",X"A6",X"7F",X"D0",X"2C",
		X"B0",X"7B",X"69",X"07",X"90",X"77",X"65",X"3F",
		X"D0",X"03",X"4C",X"79",X"16",X"69",X"FF",X"85",
		X"54",X"0A",X"65",X"54",X"A8",X"68",X"D9",X"80",
		X"02",X"B0",X"67",X"20",X"F9",X"0D",X"48",X"20",
		X"8C",X"0E",X"68",X"A4",X"7D",X"10",X"17",X"AA",
		X"F0",X"56",X"D0",X"00",X"FD",X"04",X"68",X"18",
		X"5F",X"46",X"3F",X"8A",X"2A",X"A6",X"A6",X"D0",
		X"02",X"C6",X"A7",X"C6",X"A6",X"A0",X"1B",X"85",
		X"7F",X"D0",X"D7",X"D9",X"80",X"02",X"B0",X"48",
		X"90",X"D9",X"B9",X"82",X"02",X"48",X"B9",X"81",
		X"02",X"48",X"20",X"9F",X"0E",X"A5",X"7F",X"4C",
		X"15",X"0E",X"4C",X"6E",X"0F",X"A5",X"99",X"BE",
		X"80",X"02",X"A8",X"68",X"85",X"54",X"E6",X"54",
		X"68",X"85",X"55",X"98",X"48",X"20",X"93",X"1C",
		X"A5",X"98",X"48",X"A5",X"97",X"48",X"A5",X"96",
		X"48",X"A5",X"95",X"48",X"A5",X"94",X"48",X"6C",
		X"54",X"00",X"A0",X"FF",X"68",X"F0",X"23",X"C9",
		X"64",X"F0",X"03",X"20",X"F9",X"0D",X"84",X"7D",
		X"68",X"4A",X"85",X"44",X"68",X"85",X"9C",X"68",
		X"85",X"9D",X"68",X"85",X"9E",X"68",X"85",X"9F",
		X"68",X"85",X"A0",X"68",X"85",X"A1",X"45",X"99",
		X"85",X"A2",X"A5",X"94",X"60",X"A9",X"00",X"85",
		X"3F",X"20",X"6B",X"22",X"B0",X"03",X"4C",X"6B",
		X"1D",X"20",X"5A",X"11",X"B0",X"7A",X"0F",X"00",
		X"00",X"C9",X"FF",X"D0",X"0F",X"A9",X"0E",X"A0",
		X"0F",X"20",X"1A",X"1C",X"4C",X"6B",X"22",X"82",
		X"49",X"0F",X"DA",X"A1",X"C9",X"2E",X"F0",X"E1",
		X"C9",X"A5",X"F0",X"58",X"C9",X"A4",X"F0",X"D4",
		X"C9",X"22",X"D0",X"0F",X"A5",X"A6",X"A4",X"A7",
		X"69",X"00",X"90",X"01",X"C8",X"20",X"C3",X"14",
		X"4C",X"1F",X"18",X"C9",X"A2",X"D0",X"13",X"A0",
		X"18",X"D0",X"3B",X"20",X"FD",X"11",X"A5",X"98",
		X"49",X"FF",X"A8",X"A5",X"97",X"49",X"FF",X"4C",
		X"CC",X"13",X"C9",X"9F",X"D0",X"03",X"4C",X"30",
		X"14",X"C9",X"AE",X"90",X"03",X"4C",X"EC",X"0F",
		X"20",X"60",X"0F",X"20",X"0A",X"0E",X"A9",X"29",
		X"2C",X"A9",X"28",X"2C",X"A9",X"2C",X"A0",X"00",
		X"D1",X"A6",X"D0",X"00",X"FD",X"04",X"68",X"18",
		X"03",X"4C",X"6B",X"22",X"A2",X"10",X"4C",X"4A",
		X"05",X"A0",X"15",X"68",X"68",X"4C",X"66",X"0E",
		X"20",X"D0",X"10",X"85",X"97",X"84",X"98",X"A5",
		X"77",X"A4",X"78",X"A6",X"3F",X"F0",X"21",X"A2",
		X"00",X"86",X"A3",X"C9",X"54",X"D0",X"18",X"C0",
		X"C9",X"D0",X"14",X"20",X"73",X"04",X"84",X"91",
		X"88",X"84",X"A4",X"A0",X"06",X"84",X"90",X"A0",
		X"24",X"20",X"E0",X"1E",X"4C",X"AB",X"14",X"60",
		X"A6",X"40",X"10",X"0D",X"A0",X"00",X"B1",X"97",
		X"AA",X"C8",X"B1",X"97",X"A8",X"8A",X"4C",X"CC",
		X"13",X"C9",X"54",X"D0",X"19",X"C0",X"49",X"D0",
		X"22",X"20",X"73",X"04",X"98",X"A2",X"A0",X"4C",
		X"C7",X"1C",X"A9",X"FE",X"A0",X"01",X"78",X"20",
		X"1A",X"1C",X"58",X"84",X"95",X"60",X"C9",X"53",
		X"D0",X"09",X"C0",X"54",X"D0",X"05",X"A5",X"19",
		X"4C",X"B4",X"1C",X"A5",X"97",X"A4",X"98",X"4C",
		X"1A",X"1C",X"0A",X"48",X"AA",X"20",X"6B",X"22",
		X"E0",X"83",X"90",X"20",X"20",X"60",X"0F",X"20",
		X"0A",X"0E",X"20",X"63",X"0F",X"20",X"10",X"00",
		X"00",X"FB",X"0D",X"68",X"AA",X"A5",X"98",X"48",
		X"A5",X"97",X"48",X"8A",X"48",X"20",X"DA",X"17",
		X"68",X"A8",X"8A",X"48",X"4C",X"1B",X"10",X"20",
		X"57",X"0F",X"68",X"A8",X"B9",X"F6",X"01",X"85",
		X"88",X"B9",X"F7",X"01",X"85",X"89",X"20",X"87",
		X"00",X"4C",X"F9",X"0D",X"A0",X"FF",X"2C",X"A0",
		X"00",X"84",X"3D",X"20",X"FD",X"11",X"A5",X"97",
		X"45",X"3D",X"85",X"3B",X"A5",X"98",X"45",X"3D",
		X"85",X"3C",X"20",X"74",X"1C",X"20",X"FD",X"11",
		X"A5",X"98",X"45",X"3D",X"25",X"3C",X"45",X"3D",
		X"A8",X"A5",X"97",X"45",X"3D",X"25",X"3B",X"45",
		X"3D",X"4C",X"CC",X"13",X"20",X"FC",X"0D",X"B0",
		X"13",X"A5",X"A1",X"00",X"FD",X"04",X"68",X"18",
		X"09",X"7F",X"25",X"9D",X"85",X"9D",X"A9",X"9C",
		X"A0",X"00",X"20",X"D3",X"1C",X"AA",X"4C",X"A6",
		X"10",X"A9",X"00",X"85",X"3F",X"C6",X"7F",X"20",
		X"E2",X"16",X"85",X"94",X"86",X"95",X"84",X"96",
		X"A5",X"9F",X"A4",X"A0",X"20",X"E6",X"16",X"86",
		X"9F",X"84",X"A0",X"AA",X"38",X"E5",X"94",X"F0",
		X"08",X"A9",X"01",X"90",X"04",X"A6",X"94",X"A9",
		X"FF",X"85",X"99",X"A0",X"FF",X"E8",X"C8",X"CA",
		X"D0",X"07",X"A6",X"99",X"30",X"0F",X"18",X"90",
		X"0C",X"B1",X"9F",X"D1",X"95",X"F0",X"EF",X"A2",
		X"FF",X"B0",X"02",X"A2",X"01",X"E8",X"8A",X"2A",
		X"25",X"44",X"F0",X"02",X"A9",X"FF",X"4C",X"B4",
		X"1C",X"20",X"63",X"0F",X"AA",X"20",X"D5",X"10",
		X"20",X"71",X"22",X"D0",X"F4",X"60",X"A2",X"00",
		X"20",X"71",X"22",X"86",X"3E",X"85",X"77",X"20",
		X"71",X"22",X"20",X"5A",X"11",X"B0",X"03",X"4C",
		X"6E",X"0F",X"A2",X"00",X"86",X"3F",X"86",X"40",
		X"20",X"6B",X"22",X"90",X"05",X"20",X"5A",X"11",
		X"90",X"0B",X"AA",X"20",X"6B",X"22",X"90",X"FB",
		X"20",X"5A",X"11",X"B0",X"F6",X"C9",X"11",X"00",
		X"00",X"24",X"D0",X"06",X"A9",X"FF",X"85",X"3F",
		X"D0",X"10",X"C9",X"25",X"D0",X"13",X"A5",X"42",
		X"D0",X"D0",X"A9",X"80",X"85",X"40",X"05",X"77",
		X"85",X"77",X"8A",X"09",X"80",X"AA",X"20",X"6B",
		X"22",X"86",X"78",X"38",X"05",X"42",X"E9",X"28",
		X"D0",X"03",X"4C",X"0F",X"12",X"A9",X"00",X"85",
		X"42",X"A5",X"5F",X"A6",X"60",X"A0",X"00",X"86",
		X"93",X"85",X"92",X"E4",X"62",X"D0",X"04",X"C5",
		X"61",X"F0",X"22",X"A5",X"77",X"D1",X"92",X"D0",
		X"08",X"A5",X"78",X"C8",X"D1",X"92",X"F0",X"7D",
		X"88",X"18",X"A5",X"92",X"69",X"07",X"90",X"E1",
		X"E8",X"D0",X"DC",X"00",X"FD",X"04",X"68",X"18",
		X"C9",X"41",X"90",X"05",X"E9",X"5B",X"38",X"E9",
		X"A5",X"60",X"68",X"48",X"C9",X"7C",X"D0",X"05",
		X"A9",X"8B",X"A0",X"1F",X"60",X"A5",X"77",X"A4",
		X"78",X"C9",X"54",X"D0",X"0B",X"C0",X"C9",X"F0",
		X"EF",X"C0",X"49",X"D0",X"03",X"4C",X"6E",X"0F",
		X"C9",X"53",X"D0",X"04",X"C0",X"54",X"F0",X"F5",
		X"A5",X"61",X"A4",X"62",X"85",X"92",X"84",X"93",
		X"A5",X"63",X"A4",X"64",X"85",X"8D",X"84",X"8E",
		X"18",X"69",X"07",X"90",X"01",X"C8",X"85",X"8B",
		X"84",X"8C",X"20",X"CB",X"04",X"A5",X"8B",X"A4",
		X"8C",X"C8",X"85",X"61",X"84",X"62",X"A0",X"00",
		X"A5",X"77",X"91",X"92",X"C8",X"A5",X"78",X"91",
		X"92",X"A9",X"00",X"C8",X"91",X"92",X"C8",X"91",
		X"92",X"C8",X"91",X"92",X"C8",X"91",X"92",X"C8",
		X"91",X"92",X"A5",X"92",X"18",X"69",X"02",X"A4",
		X"93",X"90",X"01",X"C8",X"85",X"79",X"84",X"7A",
		X"60",X"A5",X"3D",X"0A",X"69",X"05",X"65",X"92",
		X"A4",X"93",X"90",X"01",X"C8",X"85",X"8B",X"84",
		X"8C",X"60",X"90",X"80",X"00",X"00",X"20",X"6B",
		X"22",X"20",X"0A",X"0E",X"20",X"F9",X"0D",X"A5",
		X"99",X"30",X"0D",X"A5",X"94",X"C9",X"12",X"00",
		X"00",X"90",X"90",X"09",X"A9",X"EC",X"A0",X"11",
		X"20",X"D3",X"1C",X"D0",X"76",X"4C",X"13",X"1D",
		X"A5",X"3E",X"05",X"40",X"48",X"A5",X"3F",X"48",
		X"A0",X"00",X"98",X"48",X"A5",X"78",X"48",X"A5",
		X"77",X"48",X"20",X"F0",X"11",X"68",X"85",X"77",
		X"68",X"85",X"78",X"68",X"A8",X"BA",X"B5",X"02",
		X"48",X"B5",X"01",X"48",X"A5",X"97",X"95",X"02",
		X"A5",X"98",X"95",X"01",X"C8",X"20",X"71",X"22",
		X"C9",X"2C",X"F0",X"D6",X"84",X"3D",X"20",X"5D",
		X"0F",X"68",X"85",X"3F",X"68",X"85",X"40",X"29",
		X"7F",X"85",X"3E",X"00",X"FD",X"04",X"68",X"18",
		X"A6",X"61",X"A5",X"62",X"86",X"92",X"85",X"93",
		X"C5",X"64",X"D0",X"04",X"E4",X"63",X"F0",X"39",
		X"A0",X"00",X"B1",X"92",X"C8",X"C5",X"77",X"D0",
		X"06",X"A5",X"78",X"D1",X"92",X"F0",X"16",X"C8",
		X"B1",X"92",X"18",X"65",X"92",X"AA",X"C8",X"B1",
		X"92",X"65",X"93",X"90",X"D7",X"A2",X"6B",X"2C",
		X"A2",X"35",X"4C",X"4A",X"05",X"A2",X"78",X"A5",
		X"3E",X"D0",X"F7",X"20",X"DB",X"11",X"A5",X"3D",
		X"A0",X"04",X"D1",X"92",X"D0",X"E7",X"4C",X"25",
		X"13",X"20",X"DB",X"11",X"20",X"1B",X"05",X"A9",
		X"00",X"A8",X"85",X"A5",X"A2",X"05",X"A5",X"77",
		X"91",X"92",X"10",X"01",X"CA",X"C8",X"A5",X"78",
		X"91",X"92",X"10",X"02",X"CA",X"CA",X"86",X"A4",
		X"A5",X"3D",X"C8",X"C8",X"C8",X"91",X"92",X"A2",
		X"0B",X"A9",X"00",X"24",X"3E",X"50",X"08",X"68",
		X"18",X"69",X"01",X"AA",X"68",X"69",X"00",X"C8",
		X"91",X"92",X"C8",X"8A",X"91",X"92",X"20",X"87",
		X"13",X"86",X"A4",X"85",X"A5",X"A4",X"54",X"C6",
		X"3D",X"D0",X"DC",X"65",X"8C",X"B0",X"5D",X"85",
		X"8C",X"A8",X"8A",X"65",X"8B",X"90",X"03",X"C8",
		X"F0",X"52",X"20",X"1B",X"05",X"85",X"63",X"84",
		X"64",X"A9",X"00",X"E6",X"A5",X"A4",X"13",X"00",
		X"00",X"A4",X"F0",X"05",X"88",X"91",X"8B",X"D0",
		X"FB",X"C6",X"8C",X"C6",X"A5",X"D0",X"F5",X"E6",
		X"8C",X"38",X"A5",X"63",X"E5",X"92",X"A0",X"02",
		X"91",X"92",X"A5",X"64",X"C8",X"E5",X"93",X"91",
		X"92",X"A5",X"3E",X"D0",X"62",X"C8",X"B1",X"92",
		X"85",X"3D",X"A9",X"00",X"85",X"A4",X"85",X"A5",
		X"C8",X"68",X"AA",X"85",X"97",X"68",X"85",X"98",
		X"D1",X"92",X"90",X"0E",X"D0",X"06",X"C8",X"8A",
		X"D1",X"92",X"90",X"07",X"4C",X"7F",X"12",X"4C",
		X"48",X"05",X"C8",X"00",X"FD",X"04",X"68",X"18",
		X"A5",X"A5",X"05",X"A4",X"18",X"F0",X"0A",X"20",
		X"87",X"13",X"8A",X"65",X"97",X"AA",X"98",X"A4",
		X"54",X"65",X"98",X"86",X"A4",X"C6",X"3D",X"D0",
		X"CA",X"85",X"A5",X"A2",X"05",X"A5",X"77",X"10",
		X"01",X"CA",X"A5",X"78",X"10",X"02",X"CA",X"CA",
		X"86",X"5A",X"A9",X"00",X"20",X"90",X"13",X"8A",
		X"65",X"8B",X"85",X"79",X"98",X"65",X"8C",X"85",
		X"7A",X"A8",X"A5",X"79",X"60",X"84",X"54",X"B1",
		X"92",X"85",X"5A",X"88",X"B1",X"92",X"85",X"5B",
		X"A9",X"10",X"85",X"90",X"A2",X"00",X"A0",X"00",
		X"8A",X"0A",X"AA",X"98",X"2A",X"A8",X"B0",X"A4",
		X"06",X"A4",X"26",X"A5",X"90",X"0B",X"18",X"8A",
		X"65",X"5A",X"AA",X"98",X"65",X"5B",X"A8",X"B0",
		X"93",X"C6",X"90",X"D0",X"E3",X"60",X"A5",X"3F",
		X"F0",X"03",X"20",X"E2",X"16",X"20",X"62",X"15",
		X"38",X"A5",X"65",X"E5",X"63",X"A8",X"A5",X"66",
		X"E5",X"64",X"A2",X"00",X"86",X"3F",X"85",X"95",
		X"84",X"96",X"A2",X"90",X"4C",X"BC",X"1C",X"A5",
		X"30",X"20",X"7A",X"04",X"A9",X"00",X"F0",X"EA",
		X"A6",X"6C",X"E8",X"D0",X"9F",X"A2",X"95",X"2C",
		X"A2",X"E0",X"4C",X"4A",X"05",X"20",X"1D",X"14",
		X"20",X"E2",X"13",X"20",X"60",X"0F",X"A9",X"80",
		X"85",X"42",X"20",X"D0",X"10",X"20",X"14",X"00",
		X"00",X"F9",X"0D",X"20",X"5D",X"0F",X"A9",X"AC",
		X"20",X"65",X"0F",X"48",X"A5",X"7A",X"48",X"A5",
		X"79",X"48",X"A5",X"A7",X"48",X"A5",X"A6",X"48",
		X"20",X"E7",X"09",X"4C",X"8B",X"14",X"A9",X"9F",
		X"20",X"65",X"0F",X"09",X"80",X"85",X"42",X"20",
		X"D7",X"10",X"85",X"81",X"84",X"82",X"4C",X"F9",
		X"0D",X"20",X"1D",X"14",X"A5",X"82",X"48",X"A5",
		X"81",X"48",X"20",X"57",X"0F",X"20",X"F9",X"0D",
		X"68",X"85",X"81",X"00",X"FD",X"04",X"68",X"18",
		X"68",X"85",X"82",X"A0",X"02",X"B1",X"81",X"85",
		X"79",X"AA",X"C8",X"B1",X"81",X"F0",X"99",X"85",
		X"7A",X"C8",X"B1",X"79",X"48",X"88",X"10",X"FA",
		X"A4",X"7A",X"20",X"4C",X"1C",X"A5",X"A7",X"48",
		X"A5",X"A6",X"48",X"B1",X"81",X"85",X"A6",X"C8",
		X"B1",X"81",X"85",X"A7",X"A5",X"7A",X"48",X"A5",
		X"79",X"48",X"20",X"F6",X"0D",X"68",X"85",X"81",
		X"68",X"85",X"82",X"20",X"71",X"22",X"F0",X"03",
		X"4C",X"6E",X"0F",X"68",X"85",X"A6",X"68",X"85",
		X"A7",X"A0",X"00",X"68",X"91",X"81",X"68",X"C8",
		X"91",X"81",X"68",X"C8",X"91",X"81",X"68",X"C8",
		X"91",X"81",X"68",X"C8",X"91",X"81",X"60",X"20",
		X"F9",X"0D",X"A0",X"00",X"20",X"57",X"1E",X"68",
		X"68",X"A9",X"04",X"A0",X"02",X"D0",X"12",X"A6",
		X"97",X"A4",X"98",X"86",X"83",X"84",X"84",X"20",
		X"30",X"15",X"86",X"95",X"84",X"96",X"85",X"94",
		X"60",X"A2",X"22",X"86",X"3B",X"86",X"3C",X"85",
		X"A2",X"84",X"A3",X"85",X"95",X"84",X"96",X"A0",
		X"FF",X"C8",X"B1",X"A2",X"F0",X"0C",X"C5",X"3B",
		X"F0",X"04",X"C5",X"3C",X"D0",X"F3",X"C9",X"22",
		X"F0",X"01",X"18",X"84",X"94",X"98",X"65",X"A2",
		X"85",X"A4",X"A6",X"A3",X"90",X"01",X"E8",X"86",
		X"A5",X"A5",X"A3",X"F0",X"04",X"C9",X"24",X"D0",
		X"0B",X"98",X"20",X"B1",X"14",X"A6",X"15",X"00",
		X"00",X"A2",X"A4",X"A3",X"20",X"C4",X"16",X"A6",
		X"48",X"E0",X"54",X"D0",X"05",X"A2",X"BF",X"4C",
		X"4A",X"05",X"A5",X"94",X"95",X"00",X"A5",X"95",
		X"95",X"01",X"A5",X"96",X"95",X"02",X"A0",X"00",
		X"86",X"97",X"84",X"98",X"84",X"A3",X"88",X"84",
		X"3F",X"86",X"49",X"E8",X"E8",X"E8",X"86",X"48",
		X"60",X"46",X"41",X"48",X"49",X"FF",X"38",X"65",
		X"65",X"A4",X"66",X"00",X"FD",X"04",X"68",X"18",
		X"B0",X"01",X"88",X"C4",X"64",X"90",X"11",X"D0",
		X"04",X"C5",X"63",X"90",X"0B",X"85",X"65",X"84",
		X"66",X"85",X"67",X"84",X"68",X"AA",X"68",X"60",
		X"A2",X"4D",X"A5",X"41",X"30",X"B6",X"20",X"62",
		X"15",X"A9",X"80",X"85",X"41",X"68",X"D0",X"D0",
		X"A6",X"69",X"A5",X"6A",X"86",X"65",X"85",X"66",
		X"A0",X"00",X"84",X"82",X"84",X"81",X"A5",X"63",
		X"A6",X"64",X"85",X"92",X"86",X"93",X"A9",X"4B",
		X"A2",X"00",X"85",X"54",X"86",X"55",X"C5",X"48",
		X"F0",X"05",X"20",X"03",X"16",X"F0",X"F7",X"A9",
		X"07",X"85",X"86",X"A5",X"5F",X"A6",X"60",X"85",
		X"54",X"86",X"55",X"E4",X"62",X"D0",X"04",X"C5",
		X"61",X"F0",X"05",X"20",X"F9",X"15",X"F0",X"F3",
		X"85",X"8B",X"86",X"8C",X"A9",X"03",X"85",X"86",
		X"A5",X"8B",X"A6",X"8C",X"E4",X"64",X"D0",X"07",
		X"C5",X"63",X"D0",X"03",X"4C",X"42",X"16",X"85",
		X"54",X"86",X"55",X"A0",X"00",X"B1",X"54",X"AA",
		X"C8",X"B1",X"54",X"08",X"C8",X"B1",X"54",X"65",
		X"8B",X"85",X"8B",X"C8",X"B1",X"54",X"65",X"8C",
		X"85",X"8C",X"28",X"10",X"D3",X"8A",X"30",X"D0",
		X"C8",X"B1",X"54",X"A0",X"00",X"0A",X"69",X"05",
		X"65",X"54",X"85",X"54",X"90",X"02",X"E6",X"55",
		X"A6",X"55",X"E4",X"8C",X"D0",X"04",X"C5",X"8B",
		X"F0",X"BA",X"20",X"03",X"16",X"F0",X"F3",X"B1",
		X"54",X"30",X"35",X"C8",X"B1",X"54",X"16",X"00",
		X"00",X"10",X"30",X"C8",X"B1",X"54",X"F0",X"2B",
		X"C8",X"B1",X"54",X"AA",X"C8",X"B1",X"54",X"C5",
		X"66",X"90",X"06",X"D0",X"1E",X"E4",X"65",X"B0",
		X"1A",X"C5",X"93",X"90",X"16",X"D0",X"04",X"E4",
		X"92",X"90",X"10",X"86",X"92",X"85",X"93",X"A5",
		X"54",X"A6",X"55",X"85",X"81",X"86",X"82",X"A5",
		X"86",X"85",X"88",X"00",X"FD",X"04",X"68",X"18",
		X"A5",X"86",X"18",X"65",X"54",X"85",X"54",X"90",
		X"02",X"E6",X"55",X"A6",X"55",X"A0",X"00",X"60",
		X"A5",X"82",X"05",X"81",X"F0",X"F5",X"A5",X"88",
		X"29",X"04",X"4A",X"A8",X"85",X"88",X"B1",X"81",
		X"65",X"92",X"85",X"8D",X"A5",X"93",X"69",X"00",
		X"85",X"8E",X"A5",X"65",X"A6",X"66",X"85",X"8B",
		X"86",X"8C",X"20",X"D2",X"04",X"A4",X"88",X"C8",
		X"A5",X"8B",X"91",X"81",X"AA",X"E6",X"8C",X"A5",
		X"8C",X"C8",X"91",X"81",X"4C",X"66",X"15",X"A5",
		X"98",X"48",X"A5",X"97",X"48",X"20",X"EF",X"0E",
		X"20",X"FB",X"0D",X"68",X"85",X"A2",X"68",X"85",
		X"A3",X"A0",X"00",X"B1",X"A2",X"18",X"71",X"97",
		X"90",X"05",X"A2",X"B0",X"4C",X"4A",X"05",X"20",
		X"B1",X"14",X"20",X"B6",X"16",X"A5",X"83",X"A4",
		X"84",X"20",X"E6",X"16",X"20",X"C8",X"16",X"A5",
		X"A2",X"A4",X"A3",X"20",X"E6",X"16",X"20",X"06",
		X"15",X"4C",X"24",X"0E",X"A0",X"00",X"B1",X"A2",
		X"48",X"C8",X"B1",X"A2",X"AA",X"C8",X"B1",X"A2",
		X"A8",X"68",X"86",X"54",X"84",X"55",X"A8",X"F0",
		X"0A",X"48",X"88",X"B1",X"54",X"91",X"67",X"98",
		X"D0",X"F8",X"68",X"18",X"65",X"67",X"85",X"67",
		X"90",X"02",X"E6",X"68",X"60",X"20",X"FB",X"0D",
		X"A5",X"97",X"A4",X"98",X"85",X"54",X"84",X"55",
		X"20",X"17",X"17",X"08",X"A0",X"00",X"B1",X"54",
		X"48",X"C8",X"B1",X"54",X"AA",X"C8",X"B1",X"54",
		X"A8",X"68",X"28",X"D0",X"13",X"C4",X"17",X"00",
		X"00",X"66",X"D0",X"0F",X"E4",X"65",X"D0",X"0B",
		X"48",X"18",X"65",X"65",X"85",X"65",X"90",X"02",
		X"E6",X"66",X"68",X"86",X"54",X"84",X"55",X"60",
		X"C4",X"4A",X"D0",X"0C",X"C5",X"49",X"D0",X"08",
		X"85",X"48",X"E9",X"03",X"85",X"49",X"A0",X"00",
		X"60",X"20",X"DD",X"00",X"FD",X"04",X"68",X"18",
		X"17",X"8A",X"48",X"A9",X"01",X"20",X"B9",X"14",
		X"68",X"A0",X"00",X"91",X"95",X"68",X"68",X"4C",
		X"06",X"15",X"20",X"9D",X"17",X"D1",X"83",X"98",
		X"90",X"04",X"B1",X"83",X"AA",X"98",X"48",X"8A",
		X"48",X"20",X"B9",X"14",X"A5",X"83",X"A4",X"84",
		X"20",X"E6",X"16",X"68",X"A8",X"68",X"18",X"65",
		X"54",X"85",X"54",X"90",X"02",X"E6",X"55",X"98",
		X"20",X"C8",X"16",X"4C",X"06",X"15",X"20",X"9D",
		X"17",X"18",X"F1",X"83",X"49",X"FF",X"4C",X"42",
		X"17",X"A9",X"FF",X"85",X"98",X"20",X"71",X"22",
		X"C9",X"29",X"F0",X"06",X"20",X"63",X"0F",X"20",
		X"DA",X"17",X"20",X"9D",X"17",X"F0",X"4B",X"CA",
		X"8A",X"48",X"18",X"A2",X"00",X"F1",X"83",X"B0",
		X"B6",X"49",X"FF",X"C5",X"98",X"90",X"B1",X"A5",
		X"98",X"B0",X"AD",X"20",X"5D",X"0F",X"68",X"A8",
		X"68",X"85",X"88",X"68",X"68",X"68",X"AA",X"68",
		X"85",X"83",X"68",X"85",X"84",X"A5",X"88",X"48",
		X"98",X"48",X"A0",X"00",X"8A",X"60",X"20",X"BE",
		X"17",X"4C",X"DE",X"13",X"20",X"DF",X"16",X"A2",
		X"00",X"86",X"3F",X"A8",X"60",X"20",X"BE",X"17",
		X"F0",X"08",X"A0",X"00",X"B1",X"54",X"A8",X"4C",
		X"DE",X"13",X"4C",X"82",X"12",X"20",X"6B",X"22",
		X"20",X"F6",X"0D",X"20",X"F6",X"11",X"A6",X"97",
		X"D0",X"F0",X"A6",X"98",X"4C",X"71",X"22",X"20",
		X"BE",X"17",X"D0",X"03",X"4C",X"6F",X"19",X"A6",
		X"A6",X"A4",X"A7",X"86",X"A4",X"84",X"A5",X"A6",
		X"54",X"86",X"A6",X"18",X"65",X"54",X"18",X"00",
		X"00",X"85",X"56",X"A6",X"55",X"86",X"A7",X"90",
		X"01",X"E8",X"86",X"57",X"A0",X"00",X"B1",X"56",
		X"48",X"A9",X"00",X"91",X"56",X"20",X"71",X"22",
		X"20",X"6B",X"1D",X"68",X"A0",X"00",X"91",X"56",
		X"A6",X"A4",X"A4",X"00",X"FD",X"04",X"68",X"18",
		X"A5",X"86",X"A6",X"84",X"A7",X"60",X"20",X"F6",
		X"0D",X"20",X"34",X"18",X"20",X"63",X"0F",X"4C",
		X"DA",X"17",X"A5",X"99",X"30",X"9C",X"A5",X"94",
		X"C9",X"91",X"B0",X"96",X"20",X"13",X"1D",X"A5",
		X"97",X"A4",X"98",X"84",X"46",X"85",X"47",X"60",
		X"A5",X"47",X"48",X"A5",X"46",X"48",X"20",X"34",
		X"18",X"A0",X"00",X"EA",X"EA",X"EA",X"EA",X"EA",
		X"EA",X"EA",X"EA",X"B1",X"46",X"A8",X"68",X"85",
		X"46",X"68",X"85",X"47",X"4C",X"DE",X"13",X"20",
		X"28",X"18",X"8A",X"A0",X"00",X"91",X"46",X"60",
		X"20",X"28",X"18",X"86",X"7B",X"A2",X"00",X"20",
		X"71",X"22",X"F0",X"29",X"20",X"2E",X"18",X"86",
		X"7C",X"A0",X"00",X"B1",X"46",X"45",X"7C",X"25",
		X"7B",X"F0",X"F8",X"60",X"A9",X"89",X"A0",X"1F",
		X"4C",X"DF",X"18",X"20",X"04",X"1B",X"A5",X"99",
		X"49",X"FF",X"85",X"99",X"45",X"A1",X"85",X"A2",
		X"A5",X"94",X"4C",X"E2",X"18",X"A5",X"46",X"49",
		X"E8",X"D0",X"08",X"A2",X"14",X"45",X"47",X"49",
		X"1C",X"F0",X"0E",X"A5",X"46",X"C9",X"66",X"D0",
		X"C6",X"A5",X"47",X"E9",X"19",X"D0",X"C0",X"A2",
		X"0A",X"BD",X"E9",X"21",X"29",X"3F",X"49",X"20",
		X"18",X"69",X"20",X"20",X"00",X"2B",X"CA",X"49",
		X"21",X"D0",X"EE",X"C6",X"7B",X"D0",X"E8",X"60",
		X"20",X"11",X"1A",X"90",X"3C",X"20",X"04",X"1B",
		X"D0",X"03",X"4C",X"74",X"1C",X"A6",X"A3",X"86",
		X"89",X"A2",X"9C",X"A5",X"9C",X"A8",X"F0",X"9B",
		X"38",X"E5",X"94",X"F0",X"24",X"90",X"12",X"84",
		X"94",X"A4",X"A1",X"84",X"99",X"49",X"19",X"00",
		X"00",X"FF",X"69",X"00",X"A0",X"00",X"84",X"89",
		X"A2",X"94",X"D0",X"04",X"A0",X"00",X"84",X"A3",
		X"C9",X"F9",X"30",X"C7",X"A8",X"A5",X"A3",X"56",
		X"01",X"20",X"28",X"00",X"FD",X"04",X"68",X"18",
		X"1A",X"24",X"A2",X"10",X"57",X"A0",X"94",X"E0",
		X"9C",X"F0",X"02",X"A0",X"9C",X"38",X"49",X"FF",
		X"65",X"89",X"85",X"A3",X"B9",X"04",X"00",X"F5",
		X"04",X"85",X"98",X"B9",X"03",X"00",X"F5",X"03",
		X"85",X"97",X"B9",X"02",X"00",X"F5",X"02",X"85",
		X"96",X"B9",X"01",X"00",X"F5",X"01",X"85",X"95",
		X"B0",X"03",X"20",X"BF",X"19",X"A0",X"00",X"98",
		X"18",X"A6",X"95",X"D0",X"4A",X"A6",X"96",X"86",
		X"95",X"A6",X"97",X"86",X"96",X"A6",X"98",X"86",
		X"97",X"A6",X"A3",X"86",X"98",X"84",X"A3",X"69",
		X"08",X"C9",X"20",X"D0",X"E4",X"A9",X"00",X"85",
		X"94",X"85",X"99",X"60",X"65",X"89",X"85",X"A3",
		X"A5",X"98",X"65",X"A0",X"85",X"98",X"A5",X"97",
		X"65",X"9F",X"85",X"97",X"A5",X"96",X"65",X"9E",
		X"85",X"96",X"A5",X"95",X"65",X"9D",X"85",X"95",
		X"4C",X"AE",X"19",X"69",X"01",X"06",X"A3",X"26",
		X"98",X"26",X"97",X"26",X"96",X"26",X"95",X"10",
		X"F2",X"38",X"E5",X"94",X"B0",X"C7",X"49",X"FF",
		X"69",X"01",X"85",X"94",X"90",X"0E",X"E6",X"94",
		X"F0",X"42",X"66",X"95",X"66",X"96",X"66",X"97",
		X"66",X"98",X"66",X"A3",X"60",X"A5",X"99",X"49",
		X"FF",X"85",X"99",X"A5",X"95",X"49",X"FF",X"85",
		X"95",X"A5",X"96",X"49",X"FF",X"85",X"96",X"A5",
		X"97",X"49",X"FF",X"85",X"97",X"A5",X"98",X"49",
		X"FF",X"85",X"98",X"A5",X"A3",X"49",X"FF",X"85",
		X"A3",X"E6",X"A3",X"D0",X"0E",X"E6",X"98",X"D0",
		X"0A",X"E6",X"97",X"D0",X"06",X"E6",X"96",X"D0",
		X"02",X"E6",X"95",X"60",X"A2",X"45",X"4C",X"4A",
		X"05",X"A2",X"57",X"B4",X"04",X"84",X"1A",X"00",
		X"00",X"A3",X"B4",X"03",X"94",X"04",X"B4",X"02",
		X"94",X"03",X"B4",X"01",X"94",X"02",X"A4",X"9B",
		X"94",X"01",X"69",X"00",X"FD",X"04",X"68",X"18",
		X"08",X"30",X"E8",X"F0",X"E6",X"E9",X"08",X"A8",
		X"A5",X"A3",X"B0",X"14",X"16",X"01",X"90",X"02",
		X"F6",X"01",X"76",X"01",X"76",X"01",X"76",X"02",
		X"76",X"03",X"76",X"04",X"6A",X"C8",X"D0",X"EC",
		X"18",X"60",X"81",X"00",X"00",X"00",X"00",X"03",
		X"7F",X"5E",X"56",X"CB",X"79",X"80",X"13",X"9B",
		X"0B",X"64",X"80",X"76",X"38",X"93",X"16",X"82",
		X"38",X"AA",X"3B",X"20",X"80",X"35",X"04",X"F3",
		X"34",X"81",X"35",X"04",X"F3",X"34",X"80",X"80",
		X"00",X"00",X"00",X"80",X"31",X"72",X"17",X"F8",
		X"20",X"A3",X"1C",X"F0",X"02",X"10",X"03",X"4C",
		X"82",X"12",X"A5",X"94",X"E9",X"7F",X"48",X"A9",
		X"80",X"85",X"94",X"A9",X"4E",X"A0",X"1A",X"20",
		X"DF",X"18",X"A9",X"53",X"A0",X"1A",X"20",X"87",
		X"1B",X"A9",X"34",X"A0",X"1A",X"20",X"95",X"18",
		X"A9",X"39",X"A0",X"1A",X"20",X"99",X"20",X"A9",
		X"58",X"A0",X"1A",X"20",X"DF",X"18",X"68",X"20",
		X"F6",X"1D",X"A9",X"5D",X"A0",X"1A",X"20",X"04",
		X"1B",X"D0",X"03",X"4C",X"03",X"1B",X"20",X"2F",
		X"1B",X"A9",X"00",X"85",X"58",X"85",X"59",X"85",
		X"5A",X"85",X"5B",X"A5",X"A3",X"20",X"D1",X"1A",
		X"A5",X"98",X"20",X"D1",X"1A",X"A5",X"97",X"20",
		X"D1",X"1A",X"A5",X"96",X"20",X"D1",X"1A",X"A5",
		X"95",X"20",X"D6",X"1A",X"4C",X"07",X"1C",X"D0",
		X"03",X"4C",X"FB",X"19",X"4A",X"09",X"80",X"A8",
		X"90",X"19",X"18",X"A5",X"5B",X"65",X"A0",X"85",
		X"5B",X"A5",X"5A",X"65",X"9F",X"85",X"5A",X"A5",
		X"59",X"65",X"9E",X"85",X"59",X"A5",X"58",X"65",
		X"9D",X"85",X"58",X"66",X"58",X"66",X"59",X"66",
		X"5A",X"66",X"5B",X"66",X"A3",X"98",X"1B",X"00",
		X"00",X"4A",X"D0",X"D6",X"60",X"85",X"54",X"84",
		X"55",X"A0",X"04",X"00",X"FD",X"04",X"68",X"18",
		X"B1",X"54",X"85",X"A0",X"88",X"B1",X"54",X"85",
		X"9F",X"88",X"B1",X"54",X"85",X"9E",X"88",X"B1",
		X"54",X"85",X"A1",X"45",X"99",X"85",X"A2",X"A5",
		X"A1",X"09",X"80",X"85",X"9D",X"88",X"B1",X"54",
		X"85",X"9C",X"A5",X"94",X"60",X"A5",X"9C",X"F0",
		X"1F",X"18",X"65",X"94",X"90",X"04",X"30",X"1D",
		X"18",X"2C",X"10",X"14",X"69",X"80",X"85",X"94",
		X"D0",X"03",X"4C",X"73",X"19",X"A5",X"A2",X"85",
		X"99",X"60",X"A5",X"99",X"49",X"FF",X"30",X"05",
		X"68",X"68",X"4C",X"6F",X"19",X"4C",X"F6",X"19",
		X"20",X"84",X"1C",X"AA",X"F0",X"10",X"18",X"69",
		X"02",X"B0",X"F2",X"A2",X"00",X"86",X"A2",X"20",
		X"EF",X"18",X"E6",X"94",X"F0",X"E7",X"60",X"84",
		X"20",X"00",X"00",X"00",X"20",X"84",X"1C",X"A9",
		X"71",X"A0",X"1B",X"A2",X"00",X"86",X"A2",X"20",
		X"1A",X"1C",X"4C",X"8A",X"1B",X"20",X"04",X"1B",
		X"F0",X"76",X"20",X"93",X"1C",X"A9",X"00",X"38",
		X"E5",X"94",X"85",X"94",X"20",X"2F",X"1B",X"E6",
		X"94",X"F0",X"BA",X"A2",X"FC",X"A9",X"01",X"A4",
		X"9D",X"C4",X"95",X"D0",X"10",X"A4",X"9E",X"C4",
		X"96",X"D0",X"0A",X"A4",X"9F",X"C4",X"97",X"D0",
		X"04",X"A4",X"A0",X"C4",X"98",X"08",X"2A",X"90",
		X"09",X"E8",X"95",X"5B",X"F0",X"32",X"10",X"34",
		X"A9",X"01",X"28",X"B0",X"0E",X"06",X"A0",X"26",
		X"9F",X"26",X"9E",X"26",X"9D",X"B0",X"E6",X"30",
		X"CE",X"10",X"E2",X"A8",X"A5",X"A0",X"E5",X"98",
		X"85",X"A0",X"A5",X"9F",X"E5",X"97",X"85",X"9F",
		X"A5",X"9E",X"E5",X"96",X"85",X"9E",X"A5",X"9D",
		X"E5",X"95",X"85",X"9D",X"98",X"4C",X"C7",X"1B",
		X"A9",X"40",X"D0",X"CE",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"0A",X"85",X"A3",X"28",X"4C",X"1C",X"00",
		X"00",X"07",X"1C",X"00",X"FD",X"04",X"68",X"18",
		X"A2",X"85",X"4C",X"4A",X"05",X"A5",X"58",X"85",
		X"95",X"A5",X"59",X"85",X"96",X"A5",X"5A",X"85",
		X"97",X"A5",X"5B",X"85",X"98",X"4C",X"4F",X"19",
		X"85",X"54",X"84",X"55",X"A0",X"04",X"B1",X"54",
		X"85",X"98",X"88",X"B1",X"54",X"85",X"97",X"88",
		X"B1",X"54",X"85",X"96",X"88",X"B1",X"54",X"85",
		X"99",X"09",X"80",X"85",X"95",X"88",X"B1",X"54",
		X"85",X"94",X"84",X"A3",X"60",X"A2",X"8F",X"2C",
		X"A2",X"8A",X"A0",X"00",X"F0",X"04",X"A6",X"7B",
		X"A4",X"7C",X"20",X"93",X"1C",X"86",X"54",X"84",
		X"55",X"A0",X"04",X"A5",X"98",X"91",X"54",X"88",
		X"A5",X"97",X"91",X"54",X"88",X"A5",X"96",X"91",
		X"54",X"88",X"A5",X"99",X"09",X"7F",X"25",X"95",
		X"91",X"54",X"88",X"A5",X"94",X"91",X"54",X"84",
		X"A3",X"60",X"A5",X"A1",X"85",X"99",X"A2",X"05",
		X"B5",X"9B",X"95",X"93",X"CA",X"D0",X"F9",X"86",
		X"A3",X"60",X"20",X"93",X"1C",X"A2",X"06",X"B5",
		X"93",X"95",X"9B",X"CA",X"D0",X"F9",X"86",X"A3",
		X"60",X"A5",X"94",X"F0",X"FB",X"06",X"A3",X"90",
		X"F7",X"20",X"E7",X"19",X"D0",X"F2",X"4C",X"B0",
		X"19",X"A5",X"94",X"F0",X"09",X"A5",X"99",X"2A",
		X"A9",X"FF",X"B0",X"02",X"A9",X"01",X"60",X"20",
		X"A3",X"1C",X"85",X"95",X"A9",X"00",X"85",X"96",
		X"A2",X"88",X"A5",X"95",X"49",X"FF",X"2A",X"A9",
		X"00",X"85",X"98",X"85",X"97",X"86",X"94",X"85",
		X"A3",X"85",X"99",X"4C",X"4A",X"19",X"46",X"99",
		X"60",X"85",X"56",X"84",X"57",X"A0",X"00",X"B1",
		X"56",X"C8",X"AA",X"F0",X"C4",X"B1",X"56",X"45",
		X"99",X"30",X"C2",X"E4",X"94",X"D0",X"21",X"B1",
		X"56",X"09",X"80",X"C5",X"95",X"D0",X"19",X"C8",
		X"B1",X"56",X"C5",X"96",X"D0",X"12",X"C8",X"B1",
		X"56",X"C5",X"97",X"00",X"FD",X"04",X"68",X"18",
		X"D0",X"0B",X"C8",X"1D",X"00",X"00",X"A9",X"7F",
		X"C5",X"A3",X"B1",X"56",X"E5",X"98",X"F0",X"28",
		X"A5",X"99",X"90",X"02",X"49",X"FF",X"4C",X"A9",
		X"1C",X"A5",X"94",X"F0",X"4A",X"38",X"E9",X"A0",
		X"24",X"99",X"10",X"09",X"AA",X"A9",X"FF",X"85",
		X"9B",X"20",X"C5",X"19",X"8A",X"A2",X"94",X"C9",
		X"F9",X"10",X"06",X"20",X"11",X"1A",X"84",X"9B",
		X"60",X"A8",X"A5",X"99",X"29",X"80",X"46",X"95",
		X"05",X"95",X"85",X"95",X"20",X"28",X"1A",X"84",
		X"9B",X"60",X"A5",X"94",X"C9",X"A0",X"B0",X"20",
		X"20",X"13",X"1D",X"84",X"A3",X"A5",X"99",X"84",
		X"99",X"49",X"80",X"2A",X"A9",X"A0",X"85",X"94",
		X"A5",X"98",X"85",X"3B",X"4C",X"4A",X"19",X"85",
		X"95",X"85",X"96",X"85",X"97",X"85",X"98",X"A8",
		X"60",X"A0",X"00",X"A2",X"0A",X"94",X"90",X"CA",
		X"10",X"FB",X"90",X"0F",X"C9",X"2D",X"D0",X"04",
		X"86",X"9A",X"F0",X"04",X"C9",X"2B",X"D0",X"05",
		X"20",X"6B",X"22",X"90",X"5B",X"C9",X"2E",X"F0",
		X"2E",X"C9",X"45",X"D0",X"30",X"20",X"6B",X"22",
		X"90",X"17",X"C9",X"A5",X"F0",X"0E",X"C9",X"2D",
		X"F0",X"0A",X"C9",X"A4",X"F0",X"08",X"C9",X"2B",
		X"F0",X"04",X"D0",X"07",X"66",X"93",X"20",X"6B",
		X"22",X"90",X"5C",X"24",X"93",X"10",X"0E",X"A9",
		X"00",X"38",X"E5",X"91",X"4C",X"C1",X"1D",X"66",
		X"92",X"24",X"92",X"50",X"C3",X"A5",X"91",X"38",
		X"E5",X"90",X"85",X"91",X"F0",X"12",X"10",X"09",
		X"20",X"76",X"1B",X"E6",X"91",X"D0",X"F9",X"F0",
		X"07",X"20",X"5A",X"1B",X"C6",X"91",X"D0",X"F9",
		X"A5",X"9A",X"30",X"01",X"60",X"4C",X"0D",X"20",
		X"48",X"24",X"92",X"10",X"02",X"E6",X"90",X"20",
		X"5A",X"1B",X"68",X"38",X"E9",X"30",X"20",X"F6",
		X"1D",X"4C",X"82",X"00",X"FD",X"04",X"68",X"18",
		X"1D",X"48",X"20",X"84",X"1C",X"68",X"20",X"B4",
		X"1C",X"A5",X"A1",X"1E",X"00",X"00",X"45",X"99",
		X"85",X"A2",X"A6",X"94",X"4C",X"E2",X"18",X"A5",
		X"91",X"C9",X"0A",X"90",X"09",X"A9",X"64",X"24",
		X"93",X"30",X"11",X"4C",X"F6",X"19",X"0A",X"0A",
		X"18",X"65",X"91",X"0A",X"18",X"A0",X"00",X"71",
		X"A6",X"38",X"E9",X"30",X"85",X"91",X"4C",X"A8",
		X"1D",X"9B",X"3E",X"BC",X"1F",X"FD",X"9E",X"6E",
		X"6B",X"27",X"FD",X"9E",X"6E",X"6B",X"28",X"00",
		X"A9",X"8A",X"A0",X"04",X"20",X"52",X"1E",X"A5",
		X"6C",X"A6",X"6B",X"85",X"95",X"86",X"96",X"A2",
		X"90",X"38",X"20",X"C1",X"1C",X"20",X"55",X"1E",
		X"4C",X"EF",X"0B",X"A0",X"01",X"A9",X"20",X"24",
		X"99",X"10",X"02",X"A9",X"2D",X"99",X"04",X"02",
		X"85",X"99",X"84",X"A4",X"C8",X"A9",X"30",X"A6",
		X"94",X"D0",X"03",X"4C",X"7C",X"1F",X"A9",X"00",
		X"E0",X"80",X"F0",X"02",X"B0",X"09",X"A9",X"35",
		X"A0",X"1E",X"20",X"A0",X"1A",X"A9",X"F7",X"85",
		X"90",X"A9",X"30",X"A0",X"1E",X"20",X"D3",X"1C",
		X"F0",X"1E",X"10",X"12",X"A9",X"2B",X"A0",X"1E",
		X"20",X"D3",X"1C",X"F0",X"02",X"10",X"0E",X"20",
		X"5A",X"1B",X"C6",X"90",X"D0",X"EE",X"20",X"76",
		X"1B",X"E6",X"90",X"D0",X"DC",X"20",X"8E",X"18",
		X"20",X"13",X"1D",X"A2",X"01",X"A5",X"90",X"18",
		X"69",X"0A",X"30",X"09",X"C9",X"0B",X"B0",X"06",
		X"69",X"FF",X"AA",X"A9",X"02",X"38",X"E9",X"02",
		X"85",X"91",X"86",X"90",X"8A",X"F0",X"02",X"10",
		X"13",X"A4",X"A4",X"A9",X"2E",X"C8",X"99",X"04",
		X"02",X"8A",X"F0",X"06",X"A9",X"30",X"C8",X"99",
		X"04",X"02",X"84",X"A4",X"A0",X"00",X"A2",X"80",
		X"A5",X"98",X"18",X"79",X"91",X"1F",X"85",X"98",
		X"A5",X"97",X"79",X"00",X"FD",X"04",X"68",X"18",
		X"90",X"1F",X"85",X"97",X"A5",X"96",X"79",X"8F",
		X"1F",X"85",X"96",X"A5",X"95",X"79",X"8E",X"1F",
		X"85",X"95",X"E8",X"1F",X"00",X"00",X"B0",X"04",
		X"10",X"DE",X"30",X"02",X"30",X"DA",X"8A",X"90",
		X"04",X"49",X"FF",X"69",X"0A",X"69",X"2F",X"C8",
		X"C8",X"C8",X"C8",X"84",X"79",X"A4",X"A4",X"C8",
		X"AA",X"29",X"7F",X"99",X"04",X"02",X"C6",X"90",
		X"D0",X"06",X"A9",X"2E",X"C8",X"99",X"04",X"02",
		X"84",X"A4",X"A4",X"79",X"8A",X"49",X"FF",X"29",
		X"80",X"AA",X"C0",X"24",X"F0",X"04",X"C0",X"3C",
		X"D0",X"A6",X"A4",X"A4",X"B9",X"04",X"02",X"88",
		X"C9",X"30",X"F0",X"F8",X"C9",X"2E",X"F0",X"01",
		X"C8",X"A9",X"2B",X"A6",X"91",X"F0",X"2E",X"10",
		X"08",X"A9",X"00",X"38",X"E5",X"91",X"AA",X"A9",
		X"2D",X"99",X"06",X"02",X"A9",X"45",X"99",X"05",
		X"02",X"8A",X"A2",X"2F",X"38",X"E8",X"E9",X"0A",
		X"B0",X"FB",X"69",X"3A",X"99",X"08",X"02",X"8A",
		X"99",X"07",X"02",X"A9",X"00",X"99",X"09",X"02",
		X"F0",X"08",X"99",X"04",X"02",X"A9",X"00",X"99",
		X"05",X"02",X"A9",X"05",X"A0",X"02",X"60",X"80",
		X"00",X"00",X"00",X"00",X"FA",X"0A",X"1F",X"00",
		X"00",X"98",X"96",X"80",X"FF",X"F0",X"BD",X"C0",
		X"00",X"01",X"86",X"A0",X"FF",X"FF",X"D8",X"F0",
		X"00",X"00",X"03",X"E8",X"FF",X"FF",X"FF",X"9C",
		X"00",X"00",X"00",X"0A",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"DF",X"0A",X"80",X"00",X"03",X"4B",X"C0",
		X"FF",X"FF",X"73",X"60",X"00",X"00",X"0E",X"10",
		X"FF",X"FF",X"FD",X"A8",X"00",X"00",X"00",X"3C",
		X"20",X"84",X"1C",X"A9",X"89",X"A0",X"1F",X"20",
		X"1A",X"1C",X"F0",X"70",X"A5",X"9C",X"D0",X"03",
		X"4C",X"71",X"19",X"A2",X"81",X"A0",X"00",X"20",
		X"4C",X"1C",X"A5",X"00",X"FD",X"04",X"68",X"18",
		X"A1",X"10",X"0F",X"20",X"44",X"1D",X"A9",X"81",
		X"A0",X"00",X"20",X"D3",X"1C",X"D0",X"03",X"98",
		X"A4",X"3B",X"20",X"76",X"1C",X"98",X"48",X"20",
		X"62",X"1A",X"A9",X"20",X"00",X"00",X"81",X"A0",
		X"00",X"20",X"A0",X"1A",X"20",X"46",X"20",X"68",
		X"4A",X"90",X"0A",X"A5",X"94",X"F0",X"06",X"A5",
		X"99",X"49",X"FF",X"85",X"99",X"60",X"81",X"38",
		X"AA",X"3B",X"29",X"07",X"71",X"34",X"58",X"3E",
		X"56",X"74",X"16",X"7E",X"B3",X"1B",X"77",X"2F",
		X"EE",X"E3",X"85",X"7A",X"1D",X"84",X"1C",X"2A",
		X"7C",X"63",X"59",X"58",X"0A",X"7E",X"75",X"FD",
		X"E7",X"C6",X"80",X"31",X"72",X"18",X"10",X"81",
		X"00",X"00",X"00",X"00",X"A9",X"18",X"A0",X"20",
		X"20",X"A0",X"1A",X"A5",X"A3",X"69",X"50",X"90",
		X"03",X"20",X"9B",X"1C",X"85",X"89",X"20",X"87",
		X"1C",X"A5",X"94",X"C9",X"88",X"90",X"03",X"20",
		X"4C",X"1B",X"20",X"44",X"1D",X"A5",X"3B",X"18",
		X"69",X"81",X"F0",X"F3",X"38",X"E9",X"01",X"48",
		X"A2",X"05",X"B5",X"9C",X"B4",X"94",X"95",X"94",
		X"94",X"9C",X"CA",X"10",X"F5",X"A5",X"89",X"85",
		X"A3",X"20",X"98",X"18",X"20",X"0D",X"20",X"A9",
		X"1D",X"A0",X"20",X"20",X"AF",X"20",X"A9",X"00",
		X"85",X"A2",X"68",X"20",X"31",X"1B",X"60",X"85",
		X"A4",X"84",X"A5",X"20",X"42",X"1C",X"A9",X"8A",
		X"20",X"A0",X"1A",X"20",X"B3",X"20",X"A9",X"8A",
		X"A0",X"00",X"4C",X"A0",X"1A",X"85",X"A4",X"84",
		X"A5",X"20",X"3F",X"1C",X"B1",X"A4",X"85",X"9A",
		X"A4",X"A4",X"C8",X"98",X"D0",X"02",X"E6",X"A5",
		X"85",X"A4",X"A4",X"A5",X"20",X"A0",X"1A",X"A5",
		X"A4",X"A4",X"A5",X"18",X"69",X"05",X"90",X"01",
		X"C8",X"85",X"A4",X"84",X"A5",X"20",X"DF",X"18",
		X"A9",X"8F",X"A0",X"00",X"FD",X"04",X"68",X"18",
		X"00",X"C6",X"9A",X"D0",X"E4",X"60",X"98",X"35",
		X"44",X"7A",X"68",X"28",X"B1",X"46",X"20",X"A3",
		X"1C",X"30",X"2A",X"D0",X"13",X"A5",X"06",X"85",
		X"95",X"A5",X"0A",X"85",X"96",X"A5",X"07",X"85",
		X"97",X"A5",X"0B",X"21",X"00",X"00",X"85",X"98",
		X"4C",X"2A",X"21",X"A9",X"88",X"A0",X"22",X"20",
		X"1A",X"1C",X"A9",X"E3",X"A0",X"20",X"20",X"A0",
		X"1A",X"A9",X"E7",X"A0",X"20",X"20",X"DF",X"18",
		X"A6",X"98",X"A5",X"95",X"85",X"98",X"86",X"95",
		X"A6",X"96",X"A5",X"97",X"85",X"96",X"86",X"97",
		X"A9",X"00",X"85",X"99",X"A5",X"94",X"85",X"A3",
		X"A9",X"80",X"85",X"94",X"20",X"4F",X"19",X"A2",
		X"88",X"A0",X"22",X"4C",X"4C",X"1C",X"A9",X"BC",
		X"A0",X"21",X"20",X"DF",X"18",X"20",X"84",X"1C",
		X"A9",X"C1",X"A0",X"21",X"A6",X"A1",X"20",X"7F",
		X"1B",X"20",X"84",X"1C",X"20",X"44",X"1D",X"A9",
		X"00",X"85",X"A2",X"20",X"98",X"18",X"A9",X"C6",
		X"A0",X"21",X"20",X"95",X"18",X"A5",X"99",X"48",
		X"10",X"0D",X"20",X"8E",X"18",X"A5",X"99",X"30",
		X"09",X"A5",X"44",X"49",X"FF",X"85",X"44",X"20",
		X"0D",X"20",X"A9",X"C6",X"A0",X"21",X"20",X"DF",
		X"18",X"68",X"10",X"03",X"20",X"0D",X"20",X"A9",
		X"CB",X"A0",X"21",X"4C",X"99",X"20",X"20",X"42",
		X"1C",X"A9",X"00",X"85",X"44",X"20",X"47",X"21",
		X"A2",X"81",X"A0",X"00",X"20",X"3D",X"21",X"A9",
		X"8A",X"A0",X"00",X"20",X"1A",X"1C",X"A9",X"00",
		X"85",X"99",X"A5",X"44",X"20",X"B8",X"21",X"A9",
		X"81",X"A0",X"00",X"4C",X"87",X"1B",X"48",X"4C",
		X"79",X"21",X"81",X"49",X"0F",X"DA",X"A2",X"83",
		X"49",X"0F",X"DA",X"A2",X"7F",X"00",X"00",X"00",
		X"00",X"05",X"84",X"E6",X"1A",X"2D",X"1B",X"86",
		X"28",X"07",X"FB",X"00",X"FD",X"04",X"68",X"18",
		X"F8",X"87",X"99",X"68",X"89",X"01",X"87",X"23",
		X"35",X"DF",X"E1",X"86",X"A5",X"5D",X"E7",X"28",
		X"83",X"49",X"0F",X"DA",X"A2",X"A1",X"54",X"46",
		X"8F",X"13",X"8F",X"52",X"43",X"89",X"CD",X"E1",
		X"4E",X"8F",X"92",X"14",X"AD",X"81",X"47",X"89",
		X"C7",X"A5",X"99",X"22",X"00",X"00",X"48",X"10",
		X"03",X"20",X"0D",X"20",X"A5",X"94",X"48",X"C9",
		X"81",X"90",X"07",X"A9",X"34",X"A0",X"1A",X"20",
		X"87",X"1B",X"A9",X"2E",X"A0",X"22",X"20",X"99",
		X"20",X"68",X"C9",X"81",X"90",X"07",X"A9",X"BC",
		X"A0",X"21",X"20",X"95",X"18",X"68",X"10",X"03",
		X"4C",X"0D",X"20",X"60",X"0B",X"76",X"B3",X"83",
		X"BD",X"D3",X"79",X"1E",X"F4",X"A6",X"F5",X"7B",
		X"83",X"FC",X"B0",X"10",X"7C",X"0C",X"1F",X"67",
		X"CA",X"7C",X"DE",X"53",X"CB",X"C1",X"7D",X"14",
		X"64",X"70",X"4C",X"7D",X"B7",X"EA",X"51",X"7A",
		X"7D",X"63",X"30",X"88",X"7E",X"7E",X"92",X"44",
		X"99",X"3A",X"7E",X"4C",X"CC",X"91",X"C7",X"7F",
		X"AA",X"AA",X"AA",X"13",X"81",X"00",X"00",X"00",
		X"00",X"E6",X"A6",X"D0",X"02",X"E6",X"A7",X"84",
		X"19",X"A0",X"00",X"B1",X"A6",X"A4",X"19",X"C9",
		X"3A",X"B0",X"0A",X"C9",X"20",X"F0",X"EA",X"38",
		X"E9",X"30",X"38",X"E9",X"D0",X"60",X"80",X"4F",
		X"C7",X"52",X"58",X"A2",X"FB",X"9A",X"A9",X"4C",
		X"85",X"87",X"85",X"38",X"A9",X"82",X"A0",X"12",
		X"85",X"39",X"84",X"3A",X"A9",X"28",X"85",X"19",
		X"A9",X"1E",X"85",X"19",X"A2",X"00",X"A9",X"03",
		X"85",X"86",X"8A",X"85",X"9B",X"85",X"19",X"85",
		X"4A",X"48",X"85",X"45",X"E8",X"8E",X"02",X"24",
		X"8E",X"01",X"24",X"A2",X"4B",X"86",X"48",X"A0",
		X"71",X"85",X"5D",X"84",X"5E",X"85",X"46",X"84",
		X"47",X"A8",X"E6",X"00",X"FD",X"04",X"68",X"18",
		X"46",X"D0",X"04",X"E6",X"47",X"30",X"0F",X"A9",
		X"55",X"91",X"46",X"D1",X"46",X"D0",X"07",X"0A",
		X"91",X"46",X"D1",X"46",X"F0",X"E9",X"A5",X"01",
		X"C9",X"01",X"E9",X"00",X"85",X"47",X"A5",X"46",
		X"A4",X"47",X"85",X"69",X"84",X"6A",X"85",X"65",
		X"84",X"66",X"A2",X"00",X"A0",X"71",X"86",X"5D",
		X"84",X"5E",X"A0",X"23",X"00",X"4E",X"00",X"98",
		X"91",X"5D",X"E6",X"5D",X"A5",X"5D",X"A4",X"5E",
		X"20",X"1B",X"05",X"A9",X"3B",X"A0",X"23",X"20",
		X"EF",X"0B",X"A5",X"69",X"38",X"E5",X"5D",X"AA",
		X"A5",X"6A",X"E5",X"5E",X"20",X"45",X"1E",X"A9",
		X"2E",X"A0",X"23",X"20",X"EF",X"0B",X"20",X"44",
		X"07",X"4C",X"71",X"05",X"20",X"42",X"59",X"54",
		X"45",X"53",X"20",X"46",X"52",X"45",X"45",X"0D",
		X"00",X"23",X"23",X"23",X"20",X"4D",X"53",X"20",
		X"42",X"41",X"53",X"49",X"43",X"20",X"23",X"23",
		X"23",X"0D",X"0D",X"00",X"24",X"00",X"38",X"11",
		X"00",X"0B",X"2B",X"22",X"59",X"03",X"B4",X"E6",
		X"11",X"00",X"02",X"2B",X"30",X"59",X"00",X"F3",
		X"30",X"93",X"30",X"93",X"30",X"F3",X"30",X"11",
		X"00",X"01",X"2B",X"30",X"11",X"00",X"27",X"2B",
		X"32",X"11",X"00",X"A0",X"2B",X"24",X"11",X"60",
		X"70",X"2B",X"26",X"11",X"03",X"0B",X"2B",X"22",
		X"B4",X"F3",X"11",X"00",X"25",X"CF",X"18",X"25",
		X"00",X"54",X"11",X"00",X"01",X"2B",X"30",X"11",
		X"E0",X"01",X"2B",X"34",X"59",X"23",X"2B",X"36",
		X"21",X"34",X"35",X"50",X"1B",X"21",X"36",X"F0",
		X"30",X"93",X"36",X"21",X"34",X"90",X"23",X"59",
		X"70",X"F0",X"30",X"21",X"34",X"E3",X"10",X"E9",
		X"2B",X"34",X"93",X"30",X"93",X"30",X"1A",X"30",
		X"8C",X"F0",X"35",X"72",X"0C",X"11",X"01",X"01",
		X"2B",X"30",X"59",X"00",X"FD",X"04",X"68",X"18",
		X"60",X"F0",X"30",X"59",X"06",X"5E",X"2A",X"59",
		X"0D",X"CF",X"32",X"1A",X"2A",X"E6",X"01",X"35",
		X"4D",X"3C",X"11",X"00",X"26",X"2B",X"1A",X"11",
		X"8D",X"22",X"FF",X"26",X"00",X"47",X"2B",X"1A",
		X"11",X"0C",X"0B",X"2B",X"22",X"B4",X"E6",X"75",
		X"CF",X"32",X"63",X"90",X"00",X"11",X"E1",X"04",
		X"2B",X"22",X"11",X"00",X"0B",X"2B",X"24",X"21",
		X"30",X"2B",X"28",X"E3",X"06",X"2B",X"30",X"59",
		X"05",X"2B",X"34",X"21",X"36",X"7F",X"00",X"82",
		X"FE",X"5E",X"26",X"11",X"00",X"07",X"99",X"28",
		X"AD",X"35",X"3F",X"36",X"93",X"26",X"B4",X"CB",
		X"93",X"36",X"93",X"28",X"21",X"34",X"E6",X"01",
		X"35",X"4D",X"21",X"63",X"FF",X"27",X"00",X"59",
		X"75",X"E6",X"FF",X"35",X"3F",X"41",X"E3",X"DF",
		X"35",X"53",X"1A",X"2B",X"24",X"11",X"00",X"29",
		X"CF",X"18",X"35",X"72",X"15",X"63",X"FF",X"11",
		X"9B",X"07",X"90",X"3F",X"E6",X"5F",X"35",X"56",
		X"22",X"11",X"C0",X"FF",X"E3",X"2D",X"35",X"53",
		X"30",X"E3",X"32",X"2B",X"34",X"11",X"00",X"07",
		X"90",X"35",X"2B",X"34",X"11",X"00",X"08",X"2B",
		X"36",X"21",X"34",X"E9",X"E9",X"99",X"34",X"99",
		X"36",X"90",X"44",X"11",X"0C",X"08",X"2B",X"36",
		X"1A",X"30",X"E6",X"FB",X"35",X"56",X"52",X"11",
		X"00",X"28",X"CF",X"18",X"11",X"0F",X"26",X"CF",
		X"18",X"28",X"00",X"4C",X"11",X"E1",X"04",X"2B",
		X"22",X"11",X"00",X"0B",X"2B",X"24",X"59",X"62",
		X"5E",X"30",X"E3",X"9E",X"2B",X"34",X"AD",X"5E",
		X"31",X"21",X"30",X"E6",X"02",X"2B",X"28",X"11",
		X"00",X"07",X"99",X"28",X"AD",X"82",X"01",X"5E",
		X"26",X"B4",X"CB",X"93",X"28",X"1A",X"28",X"35",
		X"72",X"19",X"21",X"34",X"E3",X"16",X"2B",X"28",
		X"AD",X"5E",X"26",X"00",X"FD",X"04",X"68",X"18",
		X"21",X"34",X"AD",X"F0",X"28",X"1A",X"26",X"F0",
		X"34",X"93",X"34",X"93",X"34",X"1A",X"34",X"8C",
		X"DA",X"35",X"72",X"2C",X"FF",X"29",X"00",X"1F",
		X"21",X"24",X"E3",X"13",X"35",X"72",X"0D",X"75",
		X"11",X"00",X"28",X"CF",X"18",X"63",X"FF",X"E3",
		X"03",X"35",X"3F",X"1C",X"E3",X"03",X"35",X"72",
		X"1C",X"59",X"06",X"5E",X"2C",X"63",X"FF",X"2A",
		X"00",X"3E",X"A5",X"0F",X"85",X"3E",X"A5",X"0F",
		X"C5",X"3E",X"D0",X"1B",X"A5",X"0E",X"29",X"0F",
		X"D0",X"F4",X"A5",X"0E",X"29",X"10",X"D0",X"03",
		X"A9",X"20",X"2C",X"A9",X"7F",X"00",X"20",X"32",
		X"2A",X"20",X"00",X"2E",X"4C",X"04",X"2A",X"C9",
		X"FF",X"F0",X"D9",X"48",X"A9",X"20",X"00",X"20",
		X"32",X"2A",X"68",X"60",X"A5",X"30",X"38",X"E9",
		X"06",X"C9",X"60",X"90",X"02",X"85",X"30",X"60",
		X"2B",X"00",X"13",X"85",X"43",X"48",X"08",X"8A",
		X"48",X"98",X"48",X"A5",X"43",X"00",X"68",X"A8",
		X"68",X"AA",X"28",X"68",X"18",X"60",X"2C",X"00",
		X"41",X"24",X"43",X"50",X"18",X"A5",X"0F",X"C9",
		X"FF",X"69",X"00",X"C9",X"60",X"D0",X"02",X"A9",
		X"1F",X"90",X"02",X"E9",X"20",X"C9",X"0A",X"D0",
		X"02",X"A9",X"0D",X"18",X"60",X"8A",X"48",X"98",
		X"48",X"20",X"00",X"2A",X"20",X"0A",X"2C",X"C9",
		X"07",X"D0",X"04",X"00",X"4C",X"20",X"2C",X"C9",
		X"0D",X"90",X"EE",X"F0",X"03",X"48",X"00",X"68",
		X"85",X"3E",X"68",X"A8",X"68",X"AA",X"A5",X"3E",
		X"18",X"60",X"2D",X"00",X"18",X"A5",X"0F",X"C9",
		X"03",X"D0",X"03",X"4C",X"26",X"09",X"A5",X"0E",
		X"CD",X"03",X"02",X"10",X"07",X"84",X"3E",X"20",
		X"00",X"2E",X"A4",X"3E",X"60",X"2E",X"00",X"36",
		X"A5",X"0E",X"A8",X"38",X"ED",X"03",X"02",X"8C",
		X"03",X"02",X"18",X"00",X"FD",X"04",X"68",X"18",
		X"6D",X"02",X"02",X"8D",X"02",X"02",X"A9",X"00",
		X"6D",X"01",X"02",X"8D",X"01",X"02",X"A9",X"00",
		X"6D",X"00",X"02",X"8D",X"00",X"02",X"AD",X"01",
		X"02",X"C9",X"1A",X"AD",X"00",X"02",X"E9",X"4F",
		X"90",X"08",X"A9",X"00",X"8D",X"00",X"02",X"8D",
		X"01",X"02",X"60",X"2F",X"00",X"2A",X"C9",X"5F",
		X"F0",X"05",X"E0",X"5A",X"B0",X"11",X"60",X"8A",
		X"48",X"20",X"32",X"2A",X"A9",X"20",X"00",X"20",
		X"32",X"2A",X"68",X"AA",X"F0",X"08",X"CA",X"20",
		X"32",X"2A",X"90",X"03",X"A9",X"00",X"60",X"A9",
		X"3F",X"00",X"A9",X"0D",X"00",X"A2",X"00",X"60",
		X"30",X"00",X"50",X"08",X"48",X"A0",X"00",X"B9",
		X"2A",X"30",X"C8",X"20",X"00",X"2B",X"D0",X"F7",
		X"A9",X"05",X"A0",X"24",X"85",X"34",X"84",X"35",
		X"A9",X"00",X"85",X"36",X"A9",X"0A",X"85",X"37",
		X"A9",X"FE",X"A0",X"30",X"85",X"16",X"84",X"17",
		X"68",X"28",X"4C",X"9C",X"07",X"0D",X"53",X"45",
		X"4E",X"44",X"49",X"4E",X"47",X"20",X"54",X"4F",
		X"20",X"42",X"41",X"42",X"45",X"4C",X"46",X"49",
		X"53",X"48",X"0D",X"00",X"21",X"34",X"AD",X"CF",
		X"32",X"11",X"00",X"26",X"2B",X"1A",X"EE",X"00",
		X"DF",X"02",X"FF",X"31",X"00",X"5A",X"EE",X"03",
		X"F0",X"34",X"1A",X"37",X"8C",X"0A",X"35",X"72",
		X"17",X"21",X"34",X"AD",X"E6",X"20",X"35",X"56",
		X"17",X"75",X"11",X"41",X"30",X"CF",X"18",X"1A",
		X"36",X"E3",X"08",X"5E",X"36",X"21",X"34",X"AD",
		X"5E",X"37",X"93",X"34",X"8C",X"0A",X"35",X"3F",
		X"2B",X"1A",X"36",X"35",X"72",X"4F",X"11",X"05",
		X"24",X"2B",X"34",X"2B",X"24",X"59",X"01",X"5E",
		X"26",X"1A",X"36",X"5E",X"27",X"11",X"06",X"0B",
		X"2B",X"22",X"B4",X"E6",X"35",X"3F",X"4B",X"59",
		X"03",X"5E",X"0F",X"00",X"FD",X"04",X"68",X"18",
		X"59",X"00",X"5E",X"36",X"11",X"0C",X"0B",X"2B",
		X"22",X"B4",X"E6",X"90",X"FE",X"32",X"00",X"25",
		X"A0",X"00",X"B9",X"0E",X"32",X"C8",X"20",X"00",
		X"2B",X"D0",X"F7",X"4C",X"26",X"09",X"0D",X"55",
		X"53",X"45",X"20",X"42",X"41",X"42",X"45",X"4C",
		X"46",X"49",X"53",X"48",X"20",X"54",X"4F",X"20",
		X"4C",X"4F",X"41",X"44",X"00",X"00",X"00",X"4D",
		X"53",X"42",X"41",X"53",X"49",X"43",X"00",X"29",
		X"18",X"C0",X"FB",X"EE",X"19",X"02",X"00",X"C0",
		X"11",X"B4",X"26",X"2B",X"DC",X"11",X"BD",X"26",
		X"2B",X"D0",X"11",X"C6",X"26",X"2B",X"D2",X"11",
		X"CF",X"26",X"2B",X"D4",X"11",X"D8",X"26",X"2B",
		X"D6",X"11",X"E1",X"26",X"2B",X"D8",X"11",X"EA",
		X"26",X"2B",X"DA",X"11",X"20",X"0F",X"2B",X"A2",
		X"11",X"01",X"00",X"2B",X"AC",X"11",X"00",X"FF",
		X"2B",X"AE",X"11",X"00",X"00",X"2B",X"A6",X"59",
		X"00",X"5E",X"2C",X"11",X"A0",X"25",X"CF",X"18",
		X"11",X"C3",X"25",X"CF",X"18",X"59",X"00",X"2B",
		X"30",X"2B",X"32",X"2B",X"34",X"2B",X"36",X"2B",
		X"38",X"2B",X"3A",X"2B",X"3C",X"59",X"3F",X"2B",
		X"3E",X"59",X"03",X"2B",X"40",X"59",X"20",X"2B",
		X"42",X"11",X"A0",X"26",X"2B",X"84",X"59",X"3F",
		X"F3",X"84",X"11",X"A2",X"26",X"2B",X"84",X"59",
		X"2A",X"F3",X"84",X"11",X"A4",X"26",X"2B",X"84",
		X"59",X"15",X"F3",X"84",X"11",X"A6",X"26",X"2B",
		X"84",X"59",X"00",X"F3",X"84",X"11",X"AA",X"26",
		X"2B",X"84",X"59",X"03",X"F3",X"84",X"11",X"AC",
		X"26",X"2B",X"84",X"59",X"02",X"F3",X"84",X"11",
		X"AE",X"26",X"2B",X"84",X"59",X"01",X"F3",X"84",
		X"11",X"B0",X"26",X"2B",X"84",X"59",X"00",X"F3",
		X"84",X"59",X"00",X"2B",X"44",X"2B",X"46",X"59",
		X"36",X"2B",X"48",X"00",X"FD",X"04",X"68",X"18",
		X"59",X"77",X"2B",X"30",X"21",X"42",X"2B",X"B0",
		X"11",X"FF",X"FF",X"2B",X"B2",X"02",X"C0",X"37",
		X"11",X"A0",X"26",X"99",X"46",X"99",X"46",X"F6",
		X"2B",X"3E",X"11",X"AA",X"26",X"99",X"46",X"99",
		X"46",X"F6",X"2B",X"40",X"21",X"44",X"E3",X"01",
		X"2B",X"44",X"21",X"44",X"B8",X"48",X"35",X"3F",
		X"E4",X"11",X"0D",X"03",X"CF",X"18",X"21",X"46",
		X"E3",X"01",X"2B",X"46",X"59",X"00",X"2B",X"44",
		X"2B",X"DE",X"11",X"00",X"03",X"CF",X"18",X"03",
		X"00",X"0D",X"21",X"DE",X"21",X"48",X"2B",X"98",
		X"11",X"F3",X"26",X"CF",X"18",X"2B",X"48",X"03",
		X"0D",X"2C",X"21",X"30",X"2B",X"3C",X"11",X"A7",
		X"04",X"CF",X"18",X"21",X"30",X"B8",X"42",X"E3",
		X"28",X"2B",X"C0",X"11",X"90",X"01",X"2B",X"82",
		X"21",X"C0",X"2B",X"84",X"11",X"A0",X"24",X"CF",
		X"18",X"82",X"01",X"35",X"72",X"37",X"21",X"3E",
		X"FC",X"40",X"2B",X"36",X"90",X"3B",X"03",X"39",
		X"04",X"59",X"00",X"2B",X"36",X"03",X"3D",X"29",
		X"59",X"50",X"2B",X"82",X"21",X"3A",X"2B",X"84",
		X"11",X"A0",X"24",X"CF",X"18",X"21",X"92",X"2B",
		X"34",X"21",X"30",X"E3",X"08",X"2B",X"C0",X"1A",
		X"C0",X"5E",X"39",X"59",X"00",X"2B",X"32",X"21",
		X"3A",X"E3",X"9F",X"2B",X"B4",X"59",X"01",X"2B",
		X"B6",X"03",X"66",X"0D",X"21",X"34",X"35",X"72",
		X"71",X"21",X"3A",X"E6",X"01",X"2B",X"34",X"90",
		X"77",X"03",X"73",X"06",X"21",X"34",X"E6",X"01",
		X"2B",X"34",X"03",X"79",X"11",X"21",X"34",X"99",
		X"34",X"B8",X"3A",X"35",X"50",X"88",X"21",X"3E",
		X"FC",X"36",X"2B",X"4A",X"90",X"8E",X"03",X"8A",
		X"06",X"21",X"40",X"FC",X"36",X"2B",X"4A",X"03",
		X"90",X"4A",X"21",X"38",X"99",X"32",X"2B",X"C0",
		X"21",X"4A",X"F0",X"00",X"FD",X"04",X"68",X"18",
		X"C0",X"21",X"32",X"99",X"B6",X"2B",X"32",X"B8",
		X"B4",X"35",X"4D",X"A8",X"11",X"66",X"03",X"CF",
		X"18",X"21",X"30",X"99",X"30",X"2B",X"C0",X"11",
		X"F9",X"01",X"2B",X"82",X"21",X"C0",X"F0",X"82",
		X"21",X"30",X"99",X"B2",X"2B",X"30",X"B8",X"B0",
		X"35",X"50",X"C7",X"11",X"C0",X"02",X"CF",X"18",
		X"11",X"F9",X"01",X"2B",X"82",X"59",X"00",X"F0",
		X"82",X"59",X"00",X"2B",X"32",X"59",X"08",X"2B",
		X"4C",X"03",X"DA",X"1F",X"21",X"32",X"82",X"FF",
		X"2B",X"34",X"59",X"00",X"2B",X"36",X"11",X"F0",
		X"01",X"2B",X"4E",X"21",X"42",X"2B",X"3C",X"11",
		X"A7",X"04",X"CF",X"18",X"2B",X"DE",X"11",X"00",
		X"04",X"CF",X"18",X"04",X"00",X"0E",X"21",X"DE",
		X"59",X"00",X"2B",X"30",X"21",X"3A",X"2B",X"B0",
		X"59",X"01",X"2B",X"B2",X"04",X"0E",X"2E",X"21",
		X"36",X"99",X"34",X"2B",X"36",X"21",X"30",X"99",
		X"B2",X"2B",X"30",X"B8",X"B0",X"35",X"4D",X"22",
		X"11",X"0E",X"04",X"CF",X"18",X"21",X"34",X"99",
		X"34",X"2B",X"34",X"11",X"01",X"01",X"99",X"42",
		X"99",X"42",X"2B",X"4A",X"59",X"01",X"2B",X"82",
		X"11",X"A0",X"23",X"CF",X"18",X"04",X"3C",X"35",
		X"1A",X"37",X"F0",X"4A",X"21",X"36",X"82",X"FF",
		X"99",X"34",X"2B",X"36",X"21",X"4A",X"E3",X"04",
		X"2B",X"4A",X"B8",X"4E",X"35",X"53",X"56",X"11",
		X"3C",X"04",X"CF",X"18",X"59",X"11",X"AD",X"2B",
		X"82",X"59",X"00",X"2B",X"84",X"11",X"BB",X"23",
		X"CF",X"18",X"21",X"32",X"99",X"4C",X"2B",X"32",
		X"11",X"DA",X"03",X"CF",X"18",X"04",X"71",X"10",
		X"75",X"21",X"4C",X"E3",X"01",X"2B",X"4C",X"E6",
		X"20",X"35",X"56",X"7F",X"59",X"20",X"2B",X"4C",
		X"04",X"81",X"02",X"63",X"FF",X"04",X"83",X"14",
		X"75",X"21",X"4C",X"00",X"FD",X"04",X"68",X"18",
		X"E6",X"01",X"2B",X"4C",X"11",X"E0",X"FF",X"B8",
		X"4C",X"35",X"50",X"95",X"11",X"E0",X"FF",X"2B",
		X"4C",X"04",X"97",X"02",X"63",X"FF",X"04",X"99",
		X"07",X"75",X"59",X"00",X"2B",X"4C",X"63",X"FF",
		X"04",X"A0",X"07",X"75",X"59",X"00",X"2B",X"4C",
		X"63",X"FF",X"04",X"A7",X"17",X"75",X"11",X"E9",
		X"FF",X"99",X"3C",X"2B",X"3A",X"21",X"3A",X"E3",
		X"01",X"2B",X"C0",X"11",X"FE",X"FF",X"F8",X"C0",
		X"2B",X"3A",X"63",X"FF",X"04",X"BE",X"02",X"90",
		X"BC",X"22",X"A0",X"08",X"71",X"04",X"83",X"04",
		X"99",X"04",X"A0",X"04",X"22",X"A8",X"1F",X"75",
		X"59",X"08",X"2B",X"98",X"11",X"00",X"01",X"2B",
		X"9A",X"CF",X"DC",X"21",X"98",X"F3",X"9A",X"93",
		X"9A",X"93",X"9A",X"93",X"98",X"1A",X"98",X"E6",
		X"80",X"35",X"50",X"B0",X"63",X"FF",X"23",X"A0",
		X"1B",X"21",X"82",X"E6",X"01",X"2B",X"82",X"35",
		X"53",X"A8",X"FF",X"1A",X"0E",X"B8",X"AA",X"35",
		X"3F",X"A8",X"1A",X"0E",X"2B",X"AA",X"75",X"CF",
		X"DC",X"63",X"90",X"9E",X"23",X"BB",X"3A",X"75",
		X"11",X"F5",X"23",X"2B",X"86",X"2B",X"92",X"11",
		X"A0",X"22",X"2B",X"88",X"21",X"92",X"F6",X"2B",
		X"94",X"1A",X"95",X"82",X"80",X"35",X"3F",X"DB",
		X"21",X"84",X"35",X"3F",X"D9",X"CF",X"84",X"63",
		X"FF",X"21",X"94",X"B8",X"82",X"35",X"3F",X"E8",
		X"93",X"92",X"93",X"92",X"90",X"C6",X"21",X"92",
		X"B8",X"86",X"99",X"88",X"F6",X"CF",X"18",X"63",
		X"FF",X"23",X"F5",X"0A",X"FE",X"00",X"FD",X"00",
		X"BF",X"00",X"7F",X"00",X"FF",X"FF",X"24",X"A0",
		X"5A",X"21",X"82",X"FC",X"84",X"2B",X"94",X"21",
		X"82",X"35",X"53",X"AF",X"59",X"00",X"B8",X"82",
		X"2B",X"82",X"21",X"84",X"35",X"53",X"BA",X"59",
		X"00",X"B8",X"84",X"00",X"FD",X"04",X"68",X"18",
		X"2B",X"84",X"59",X"00",X"2B",X"92",X"2B",X"96",
		X"21",X"92",X"99",X"92",X"2B",X"92",X"21",X"82",
		X"35",X"53",X"CD",X"93",X"92",X"21",X"82",X"99",
		X"82",X"2B",X"82",X"21",X"92",X"B8",X"84",X"35",
		X"50",X"DE",X"2B",X"92",X"93",X"82",X"75",X"CF",
		X"DC",X"63",X"21",X"96",X"E3",X"01",X"82",X"0F",
		X"35",X"72",X"BE",X"21",X"94",X"35",X"53",X"F5",
		X"59",X"00",X"B8",X"82",X"FF",X"21",X"82",X"FF",
		X"25",X"A0",X"23",X"75",X"11",X"A8",X"22",X"CF",
		X"18",X"11",X"02",X"00",X"2B",X"A4",X"11",X"FF",
		X"7F",X"F8",X"AC",X"2B",X"AC",X"1A",X"A2",X"5E",
		X"24",X"5E",X"25",X"5E",X"26",X"5E",X"27",X"11",
		X"D4",X"04",X"2B",X"22",X"63",X"FF",X"25",X"C3",
		X"3A",X"75",X"11",X"A0",X"25",X"CF",X"18",X"11",
		X"00",X"08",X"2B",X"28",X"1A",X"29",X"5E",X"94",
		X"CF",X"DC",X"1A",X"94",X"5E",X"29",X"B4",X"FF",
		X"11",X"87",X"00",X"B8",X"94",X"5E",X"29",X"B4",
		X"FF",X"1A",X"28",X"E3",X"04",X"5E",X"28",X"E6",
		X"A0",X"35",X"50",X"D0",X"59",X"00",X"5E",X"28",
		X"93",X"94",X"1A",X"94",X"E6",X"44",X"35",X"50",
		X"D0",X"63",X"FF",X"26",X"A0",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"26",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"26",X"B4",X"09",
		X"75",X"11",X"BC",X"26",X"CF",X"18",X"63",X"FF",
		X"FF",X"26",X"BD",X"09",X"35",X"3F",X"C1",X"59",
		X"00",X"FF",X"59",X"01",X"FF",X"26",X"C6",X"09",
		X"35",X"72",X"CA",X"59",X"00",X"FF",X"59",X"01",
		X"FF",X"26",X"CF",X"09",X"35",X"56",X"D3",X"59",
		X"00",X"FF",X"59",X"01",X"FF",X"26",X"D8",X"09",
		X"35",X"53",X"DC",X"59",X"00",X"FF",X"59",X"01",
		X"FF",X"26",X"E1",X"00",X"FD",X"04",X"68",X"18",
		X"09",X"35",X"50",X"E5",X"59",X"00",X"FF",X"59",
		X"01",X"FF",X"26",X"EA",X"09",X"35",X"4D",X"EE",
		X"59",X"00",X"FF",X"59",X"01",X"FF",X"26",X"F3",
		X"0A",X"11",X"00",X"06",X"2B",X"22",X"21",X"98",
		X"B4",X"F6",X"FF",X"00",X"00",X"45",X"67",X"67",
		X"00",X"00",X"00",X"00",X"00",X"45",X"18",X"E6",
		X"FB",X"EE",X"19",X"02",X"00",X"18",X"1A",X"21",
		X"E6",X"F8",X"35",X"53",X"0B",X"21",X"0E",X"F3",
		X"17",X"90",X"05",X"11",X"00",X"05",X"2B",X"30",
		X"11",X"A0",X"58",X"2B",X"1A",X"FF",X"58",X"A0",
		X"38",X"CD",X"D1",X"75",X"CD",X"AA",X"43",X"4D",
		X"44",X"30",X"20",X"20",X"00",X"CF",X"32",X"59",
		X"00",X"2B",X"34",X"59",X"0A",X"2B",X"36",X"CF",
		X"38",X"21",X"36",X"E6",X"01",X"35",X"4D",X"B2",
		X"CF",X"3A",X"CD",X"C7",X"40",X"00",X"00",X"00",
		X"00",X"95",X"CF",X"3C",X"CF",X"3E",X"8C",X"01",
		X"CF",X"40",X"63",X"FF",X"2B",X"42",X"93",X"1B",
		X"FF",X"59",X"A0",X"4C",X"CD",X"E5",X"75",X"CD",
		X"AA",X"43",X"4D",X"44",X"38",X"20",X"20",X"00",
		X"CF",X"32",X"CF",X"3A",X"CD",X"B6",X"48",X"00",
		X"00",X"01",X"AA",X"87",X"CF",X"3C",X"CF",X"3E",
		X"8C",X"FF",X"35",X"3F",X"DD",X"21",X"44",X"82",
		X"04",X"35",X"3F",X"CC",X"59",X"01",X"2B",X"34",
		X"90",X"DD",X"CF",X"38",X"CF",X"38",X"CF",X"38",
		X"CF",X"38",X"8C",X"AA",X"35",X"72",X"DD",X"59",
		X"02",X"2B",X"34",X"21",X"44",X"82",X"FA",X"CF",
		X"40",X"63",X"FF",X"2B",X"46",X"93",X"1B",X"FF",
		X"5A",X"A0",X"5C",X"CD",X"D3",X"75",X"CD",X"AA",
		X"43",X"4D",X"44",X"35",X"38",X"20",X"00",X"CF",
		X"32",X"CF",X"3A",X"CD",X"B6",X"7A",X"00",X"00",
		X"00",X"00",X"00",X"CF",X"3C",X"CF",X"3E",X"CF",
		X"38",X"CF",X"38",X"00",X"FD",X"04",X"68",X"18",
		X"CF",X"38",X"82",X"C0",X"8C",X"C0",X"35",X"72",
		X"CB",X"59",X"04",X"2B",X"34",X"21",X"44",X"82",
		X"FE",X"CF",X"40",X"63",X"FF",X"2B",X"48",X"CD",
		X"F5",X"75",X"CD",X"E1",X"43",X"4D",X"44",X"35",
		X"35",X"20",X"00",X"CF",X"32",X"CD",X"EB",X"77",
		X"00",X"00",X"00",X"00",X"00",X"CF",X"3C",X"CF",
		X"3E",X"82",X"FE",X"CF",X"40",X"63",X"FF",X"2B",
		X"4A",X"93",X"1B",X"FF",X"5B",X"A0",X"58",X"CD",
		X"CF",X"75",X"CD",X"AA",X"41",X"43",X"4D",X"44",
		X"34",X"31",X"00",X"CF",X"32",X"21",X"34",X"8C",
		X"01",X"35",X"72",X"BD",X"CD",X"BB",X"69",X"00",
		X"00",X"00",X"00",X"00",X"90",X"C5",X"CD",X"C5",
		X"69",X"40",X"00",X"00",X"00",X"00",X"CF",X"3C",
		X"CF",X"3E",X"82",X"FE",X"CF",X"40",X"63",X"FF",
		X"2B",X"4C",X"CD",X"F1",X"75",X"CD",X"DD",X"43",
		X"4D",X"44",X"31",X"36",X"20",X"00",X"CF",X"32",
		X"CD",X"E7",X"50",X"00",X"00",X"02",X"00",X"00",
		X"CF",X"3C",X"CF",X"3E",X"82",X"FE",X"CF",X"40",
		X"63",X"FF",X"2B",X"4E",X"93",X"1B",X"FF",X"5C",
		X"A0",X"40",X"CD",X"D9",X"75",X"CD",X"A9",X"51",
		X"00",X"00",X"00",X"00",X"00",X"2B",X"50",X"2B",
		X"52",X"1A",X"55",X"93",X"52",X"F0",X"52",X"1A",
		X"54",X"93",X"52",X"F0",X"52",X"1A",X"57",X"93",
		X"52",X"F0",X"52",X"1A",X"56",X"93",X"52",X"F0",
		X"52",X"21",X"50",X"CF",X"3C",X"CF",X"3E",X"82",
		X"FE",X"35",X"72",X"D7",X"CF",X"38",X"8C",X"FF",
		X"35",X"3F",X"D0",X"63",X"FF",X"2B",X"58",X"93",
		X"1B",X"FF",X"5D",X"A0",X"3B",X"CD",X"AB",X"11",
		X"09",X"0B",X"2B",X"22",X"11",X"78",X"80",X"B4",
		X"FA",X"FF",X"2B",X"3A",X"CD",X"BA",X"11",X"09",
		X"0B",X"2B",X"22",X"11",X"7C",X"80",X"B4",X"FA",
		X"FF",X"2B",X"5A",X"00",X"FD",X"04",X"68",X"18",
		X"CD",X"D4",X"59",X"FF",X"5E",X"2A",X"59",X"2A",
		X"2B",X"24",X"E3",X"01",X"2B",X"26",X"11",X"15",
		X"0B",X"2B",X"22",X"B4",X"CB",X"1A",X"2A",X"FF",
		X"2B",X"38",X"93",X"1B",X"FF",X"5E",X"A0",X"2B",
		X"CD",X"C4",X"FC",X"5D",X"5E",X"5D",X"59",X"08",
		X"2B",X"36",X"21",X"5C",X"35",X"53",X"B8",X"99",
		X"5C",X"2B",X"5C",X"11",X"21",X"10",X"FC",X"5C",
		X"90",X"BA",X"99",X"5C",X"2B",X"5C",X"21",X"36",
		X"E6",X"01",X"35",X"4D",X"A6",X"FF",X"2B",X"5E",
		X"93",X"1B",X"FF",X"5F",X"A0",X"5E",X"CD",X"D6",
		X"75",X"2B",X"50",X"21",X"60",X"2B",X"52",X"59",
		X"FF",X"F0",X"52",X"93",X"52",X"F0",X"52",X"93",
		X"52",X"59",X"06",X"2B",X"36",X"21",X"50",X"AD",
		X"93",X"50",X"F0",X"52",X"93",X"52",X"21",X"36",
		X"E6",X"01",X"35",X"4D",X"B3",X"21",X"60",X"2B",
		X"24",X"E3",X"08",X"2B",X"26",X"11",X"15",X"0B",
		X"2B",X"22",X"B4",X"CB",X"63",X"FF",X"2B",X"3C",
		X"CD",X"F7",X"75",X"59",X"08",X"2B",X"36",X"CF",
		X"38",X"82",X"80",X"35",X"3F",X"ED",X"21",X"36",
		X"E6",X"01",X"35",X"4D",X"DD",X"1A",X"2A",X"2B",
		X"44",X"CF",X"62",X"21",X"44",X"63",X"FF",X"2B",
		X"3E",X"93",X"1B",X"FF",X"60",X"A0",X"5C",X"CD",
		X"D0",X"75",X"CF",X"42",X"35",X"3F",X"AF",X"CF",
		X"5A",X"1A",X"0E",X"E6",X"3C",X"35",X"50",X"A1",
		X"CF",X"46",X"CF",X"4A",X"CF",X"4C",X"21",X"44",
		X"35",X"3F",X"C1",X"1A",X"0E",X"E6",X"78",X"35",
		X"50",X"B1",X"21",X"34",X"8C",X"02",X"35",X"72",
		X"CA",X"CF",X"48",X"CF",X"4E",X"CF",X"5A",X"63",
		X"FF",X"2B",X"64",X"CD",X"F5",X"75",X"CF",X"66",
		X"CD",X"E1",X"56",X"6F",X"6C",X"2E",X"49",X"44",
		X"20",X"00",X"CF",X"32",X"59",X"0B",X"99",X"30",
		X"F6",X"2B",X"68",X"00",X"FD",X"04",X"68",X"18",
		X"CF",X"6A",X"11",X"00",X"02",X"FC",X"68",X"CF",
		X"40",X"63",X"FF",X"2B",X"6C",X"93",X"1B",X"FF",
		X"61",X"A0",X"4E",X"CD",X"E7",X"75",X"59",X"00",
		X"2B",X"56",X"2B",X"54",X"CF",X"66",X"CD",X"B0",
		X"4D",X"42",X"52",X"20",X"00",X"CF",X"32",X"11",
		X"FE",X"01",X"99",X"30",X"F6",X"2B",X"68",X"11",
		X"55",X"AA",X"FC",X"68",X"35",X"72",X"E5",X"11",
		X"C6",X"01",X"99",X"30",X"F6",X"2B",X"56",X"11",
		X"C8",X"01",X"99",X"30",X"F6",X"2B",X"54",X"11",
		X"C2",X"01",X"99",X"30",X"AD",X"2B",X"68",X"CF",
		X"62",X"59",X"0B",X"FC",X"68",X"35",X"3F",X"E5",
		X"8C",X"07",X"63",X"FF",X"2B",X"6E",X"93",X"1B",
		X"FF",X"62",X"A0",X"5F",X"CD",X"FA",X"75",X"59",
		X"0D",X"99",X"30",X"AD",X"2B",X"70",X"21",X"56",
		X"2B",X"72",X"21",X"54",X"2B",X"74",X"59",X"0E",
		X"99",X"30",X"F6",X"2B",X"76",X"59",X"00",X"2B",
		X"78",X"CF",X"7A",X"2B",X"7C",X"21",X"74",X"2B",
		X"7E",X"59",X"24",X"99",X"30",X"F6",X"2B",X"76",
		X"59",X"26",X"99",X"30",X"F6",X"2B",X"78",X"CF",
		X"7A",X"CF",X"7A",X"59",X"00",X"B8",X"70",X"B8",
		X"70",X"2B",X"76",X"11",X"FF",X"FF",X"2B",X"78",
		X"CF",X"7A",X"2B",X"81",X"21",X"74",X"2B",X"83",
		X"59",X"2C",X"99",X"30",X"F6",X"2B",X"85",X"59",
		X"2E",X"99",X"30",X"F6",X"2B",X"87",X"63",X"FF",
		X"93",X"1B",X"FF",X"63",X"A0",X"52",X"2B",X"89",
		X"CD",X"B6",X"75",X"CF",X"3A",X"21",X"34",X"E6",
		X"02",X"35",X"53",X"AE",X"CF",X"8B",X"CF",X"58",
		X"59",X"00",X"2B",X"5C",X"63",X"FF",X"2B",X"8D",
		X"CD",X"EB",X"75",X"CF",X"8D",X"21",X"30",X"2B",
		X"52",X"59",X"00",X"2B",X"5C",X"11",X"00",X"02",
		X"2B",X"68",X"CF",X"38",X"F0",X"52",X"CF",X"5E",
		X"21",X"52",X"E3",X"00",X"FD",X"04",X"68",X"18",
		X"01",X"2B",X"52",X"21",X"68",X"E6",X"01",X"35",
		X"4D",X"C8",X"CF",X"38",X"CF",X"5E",X"CF",X"38",
		X"CF",X"5E",X"CF",X"5A",X"21",X"5C",X"63",X"FF",
		X"2B",X"66",X"93",X"1B",X"FF",X"64",X"A0",X"52",
		X"CD",X"D6",X"75",X"21",X"8F",X"FC",X"91",X"35",
		X"72",X"AC",X"21",X"93",X"FC",X"95",X"35",X"3F",
		X"D2",X"11",X"FF",X"01",X"F8",X"8F",X"35",X"72",
		X"BF",X"CF",X"38",X"CF",X"38",X"CF",X"8D",X"CF",
		X"97",X"21",X"8F",X"E3",X"01",X"2B",X"8F",X"35",
		X"72",X"CE",X"21",X"93",X"E3",X"01",X"2B",X"93",
		X"CF",X"38",X"90",X"D4",X"E6",X"01",X"63",X"FF",
		X"2B",X"99",X"CD",X"EB",X"75",X"21",X"85",X"2B",
		X"72",X"21",X"87",X"2B",X"74",X"CF",X"9B",X"CF",
		X"66",X"93",X"56",X"63",X"FF",X"2B",X"9D",X"93",
		X"1B",X"FF",X"65",X"A0",X"60",X"CD",X"C9",X"75",
		X"59",X"00",X"2B",X"8F",X"2B",X"93",X"21",X"50",
		X"E3",X"1C",X"F6",X"2B",X"91",X"21",X"50",X"E3",
		X"1E",X"F6",X"2B",X"95",X"21",X"50",X"E3",X"1A",
		X"F6",X"2B",X"72",X"21",X"50",X"E3",X"14",X"F6",
		X"2B",X"74",X"CF",X"9F",X"CF",X"9B",X"63",X"FF",
		X"2B",X"A1",X"CD",X"F9",X"75",X"1A",X"75",X"82",
		X"0F",X"5E",X"75",X"59",X"01",X"2B",X"68",X"B8",
		X"70",X"35",X"53",X"E5",X"CF",X"A3",X"21",X"68",
		X"99",X"68",X"90",X"D6",X"21",X"81",X"2B",X"76",
		X"21",X"83",X"2B",X"78",X"CF",X"7A",X"21",X"72",
		X"2B",X"56",X"21",X"74",X"2B",X"54",X"63",X"FF",
		X"2B",X"9B",X"93",X"1B",X"FF",X"66",X"A0",X"5F",
		X"CD",X"BD",X"75",X"59",X"00",X"5E",X"76",X"1A",
		X"72",X"5E",X"77",X"1A",X"73",X"5E",X"78",X"1A",
		X"74",X"5E",X"79",X"21",X"76",X"2B",X"72",X"21",
		X"78",X"2B",X"74",X"CF",X"7A",X"63",X"FF",X"2B",
		X"8B",X"CD",X"D0",X"00",X"FD",X"04",X"68",X"18",
		X"75",X"21",X"72",X"2B",X"76",X"21",X"74",X"2B",
		X"78",X"CF",X"7A",X"21",X"78",X"63",X"FF",X"2B",
		X"A3",X"CD",X"FA",X"21",X"72",X"FC",X"76",X"35",
		X"53",X"DF",X"21",X"72",X"90",X"E2",X"11",X"00",
		X"80",X"99",X"76",X"35",X"50",X"ED",X"21",X"74",
		X"E3",X"01",X"2B",X"74",X"21",X"74",X"99",X"78",
		X"2B",X"74",X"21",X"72",X"99",X"76",X"2B",X"72",
		X"FF",X"93",X"1B",X"FF",X"67",X"A0",X"42",X"2B",
		X"7A",X"CD",X"B9",X"75",X"E6",X"20",X"35",X"53",
		X"AC",X"59",X"7F",X"90",X"B3",X"E6",X"60",X"35",
		X"50",X"B3",X"59",X"7F",X"82",X"7F",X"CF",X"A5",
		X"63",X"FF",X"2B",X"A7",X"CD",X"CA",X"75",X"21",
		X"74",X"CF",X"6A",X"21",X"72",X"CF",X"6A",X"CF",
		X"A9",X"63",X"FF",X"2B",X"AB",X"CD",X"DB",X"75",
		X"2B",X"68",X"1A",X"69",X"CF",X"62",X"1A",X"68",
		X"CF",X"62",X"63",X"FF",X"2B",X"6A",X"93",X"1B",
		X"FF",X"68",X"A0",X"56",X"CD",X"B5",X"75",X"DF",
		X"FE",X"EC",X"00",X"E9",X"E9",X"E9",X"E9",X"1A",
		X"19",X"CF",X"AD",X"EE",X"00",X"DF",X"02",X"CF",
		X"AD",X"63",X"FF",X"2B",X"62",X"CD",X"D9",X"75",
		X"2B",X"68",X"35",X"72",X"C8",X"CD",X"C6",X"20",
		X"4F",X"4B",X"0A",X"00",X"90",X"D3",X"CD",X"D3",
		X"20",X"46",X"41",X"49",X"4C",X"45",X"44",X"0A",
		X"00",X"CF",X"32",X"21",X"68",X"63",X"FF",X"2B",
		X"40",X"CD",X"EF",X"75",X"82",X"0F",X"E6",X"0A",
		X"35",X"53",X"E9",X"E3",X"3A",X"90",X"EB",X"E3",
		X"41",X"CF",X"A5",X"63",X"FF",X"2B",X"AD",X"93",
		X"1B",X"FF",X"69",X"A0",X"4E",X"CD",X"BC",X"75",
		X"2B",X"52",X"21",X"52",X"AD",X"35",X"3F",X"BA",
		X"8C",X"0A",X"35",X"3F",X"B4",X"8C",X"0A",X"CF",
		X"A5",X"90",X"B6",X"CF",X"A9",X"93",X"52",X"90",
		X"A3",X"63",X"FF",X"00",X"FD",X"04",X"68",X"18",
		X"2B",X"32",X"CD",X"E7",X"75",X"CD",X"CB",X"56",
		X"6F",X"6C",X"75",X"6D",X"65",X"20",X"00",X"CF",
		X"32",X"21",X"50",X"2B",X"52",X"59",X"0B",X"2B",
		X"68",X"21",X"52",X"AD",X"93",X"52",X"CF",X"A7",
		X"21",X"68",X"E6",X"01",X"35",X"4D",X"D3",X"CF",
		X"A9",X"63",X"FF",X"2B",X"AF",X"93",X"1B",X"FF",
		X"6A",X"A0",X"4F",X"CD",X"B3",X"75",X"2B",X"B1",
		X"59",X"30",X"2B",X"68",X"59",X"0A",X"CF",X"B3",
		X"21",X"B1",X"E3",X"30",X"CF",X"A5",X"63",X"FF",
		X"2B",X"B5",X"CD",X"E8",X"75",X"11",X"00",X"06",
		X"2B",X"22",X"21",X"50",X"E3",X"11",X"AD",X"B4",
		X"F6",X"E6",X"14",X"35",X"53",X"CB",X"E3",X"64",
		X"CF",X"B5",X"11",X"6D",X"06",X"2B",X"22",X"21",
		X"50",X"E3",X"10",X"F6",X"B4",X"F5",X"82",X"0F",
		X"CF",X"B5",X"21",X"50",X"E3",X"10",X"AD",X"82",
		X"1F",X"CF",X"B5",X"63",X"FF",X"2B",X"B7",X"93",
		X"1B",X"FF",X"6B",X"A0",X"53",X"CD",X"B7",X"75",
		X"CF",X"B7",X"59",X"04",X"99",X"B9",X"2B",X"B9",
		X"CF",X"BB",X"59",X"04",X"99",X"B9",X"2B",X"B9",
		X"CF",X"BD",X"CF",X"A9",X"63",X"FF",X"2B",X"BF",
		X"CD",X"EC",X"75",X"21",X"50",X"2B",X"52",X"59",
		X"0B",X"2B",X"68",X"8C",X"03",X"35",X"72",X"D5",
		X"21",X"52",X"AD",X"8C",X"20",X"35",X"3F",X"D5",
		X"59",X"2E",X"CF",X"A5",X"21",X"52",X"AD",X"93",
		X"52",X"8C",X"20",X"35",X"3F",X"E3",X"8C",X"20",
		X"CF",X"A7",X"21",X"68",X"E6",X"01",X"35",X"4D",
		X"C2",X"63",X"FF",X"2B",X"BD",X"93",X"1B",X"FF",
		X"6C",X"A0",X"2C",X"CD",X"C5",X"75",X"2B",X"36",
		X"21",X"B1",X"B8",X"36",X"35",X"50",X"B0",X"2B",
		X"B1",X"93",X"68",X"90",X"A5",X"21",X"68",X"35",
		X"72",X"BB",X"59",X"20",X"CF",X"A5",X"90",X"C3",
		X"88",X"30",X"CF",X"00",X"FD",X"04",X"68",X"18",
		X"A5",X"59",X"30",X"2B",X"68",X"63",X"FF",X"2B",
		X"B3",X"93",X"1B",X"FF",X"6D",X"A0",X"4E",X"CD",
		X"E7",X"11",X"20",X"3F",X"2B",X"24",X"59",X"00",
		X"5E",X"B9",X"11",X"20",X"01",X"AD",X"5E",X"BA",
		X"21",X"B9",X"2B",X"28",X"5E",X"26",X"11",X"E1",
		X"04",X"2B",X"22",X"B4",X"CB",X"93",X"28",X"1A",
		X"28",X"8C",X"A0",X"35",X"72",X"B5",X"59",X"01",
		X"5E",X"37",X"59",X"D0",X"E3",X"1E",X"5E",X"36",
		X"21",X"36",X"AD",X"E6",X"78",X"35",X"53",X"DB",
		X"E3",X"80",X"90",X"DD",X"E3",X"18",X"F0",X"36",
		X"1A",X"36",X"E6",X"20",X"35",X"4D",X"CB",X"FF",
		X"2B",X"A9",X"93",X"1B",X"FF",X"6E",X"A0",X"50",
		X"CD",X"E9",X"E6",X"52",X"35",X"53",X"AE",X"E3",
		X"32",X"2B",X"36",X"11",X"00",X"07",X"90",X"B3",
		X"2B",X"36",X"11",X"00",X"08",X"2B",X"C1",X"21",
		X"36",X"E9",X"E9",X"99",X"36",X"99",X"C1",X"2B",
		X"C1",X"11",X"20",X"3F",X"2B",X"24",X"21",X"B9",
		X"2B",X"28",X"E3",X"06",X"2B",X"B9",X"11",X"E1",
		X"04",X"2B",X"22",X"59",X"05",X"2B",X"36",X"21",
		X"C1",X"7F",X"00",X"5E",X"26",X"B4",X"CB",X"93",
		X"C1",X"93",X"28",X"21",X"36",X"E6",X"01",X"35",
		X"4D",X"D3",X"FF",X"2B",X"A5",X"93",X"1B",X"FF",
		X"6F",X"A0",X"58",X"CD",X"F1",X"75",X"21",X"30",
		X"2B",X"50",X"11",X"00",X"02",X"99",X"30",X"B8",
		X"50",X"35",X"4D",X"B7",X"CF",X"66",X"93",X"56",
		X"21",X"30",X"90",X"A3",X"21",X"50",X"AD",X"35",
		X"3F",X"EF",X"8C",X"E5",X"35",X"3F",X"E9",X"21",
		X"50",X"E3",X"0B",X"AD",X"2B",X"68",X"8C",X"0F",
		X"35",X"3F",X"E9",X"82",X"02",X"35",X"3F",X"E9",
		X"21",X"68",X"82",X"08",X"35",X"3F",X"DE",X"CF",
		X"AF",X"90",X"E9",X"CF",X"BF",X"CF",X"C3",X"35",
		X"72",X"E9",X"CF",X"00",X"FD",X"04",X"68",X"18",
		X"C5",X"CF",X"C7",X"21",X"50",X"E3",X"20",X"90",
		X"A3",X"63",X"FF",X"2B",X"C9",X"93",X"1B",X"FF",
		X"70",X"A0",X"5E",X"CD",X"F7",X"75",X"21",X"50",
		X"E3",X"0B",X"AD",X"82",X"10",X"35",X"3F",X"B7",
		X"CD",X"B5",X"20",X"20",X"3C",X"44",X"49",X"52",
		X"3E",X"00",X"90",X"F3",X"21",X"50",X"E3",X"1C",
		X"F6",X"2B",X"72",X"21",X"50",X"E3",X"1E",X"F6",
		X"2B",X"74",X"CF",X"CB",X"59",X"00",X"2B",X"C1",
		X"59",X"08",X"2B",X"36",X"21",X"52",X"AD",X"8C",
		X"30",X"35",X"72",X"EF",X"21",X"36",X"E6",X"06",
		X"35",X"53",X"E4",X"59",X"20",X"F0",X"52",X"90",
		X"E6",X"93",X"C1",X"93",X"52",X"21",X"36",X"E6",
		X"01",X"35",X"53",X"CD",X"21",X"60",X"99",X"C1",
		X"CF",X"32",X"63",X"FF",X"2B",X"BB",X"93",X"1B",
		X"FF",X"71",X"A0",X"5F",X"CD",X"FA",X"75",X"59",
		X"09",X"2B",X"36",X"21",X"60",X"99",X"36",X"2B",
		X"52",X"59",X"30",X"F0",X"52",X"21",X"36",X"E6",
		X"01",X"35",X"53",X"A3",X"59",X"1F",X"2B",X"C1",
		X"CF",X"A3",X"35",X"50",X"C3",X"59",X"6A",X"90",
		X"C5",X"59",X"69",X"2B",X"68",X"59",X"09",X"2B",
		X"36",X"21",X"60",X"99",X"36",X"2B",X"52",X"21",
		X"52",X"AD",X"E9",X"B8",X"68",X"35",X"53",X"E2",
		X"E3",X"3A",X"F0",X"52",X"59",X"6A",X"90",X"E8",
		X"E3",X"30",X"F0",X"52",X"59",X"69",X"2B",X"68",
		X"21",X"36",X"E6",X"01",X"35",X"53",X"C9",X"21",
		X"C1",X"E6",X"01",X"35",X"53",X"B8",X"63",X"FF",
		X"93",X"1B",X"FF",X"72",X"A0",X"14",X"2B",X"CB",
		X"CD",X"AD",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",
		X"2D",X"2D",X"2D",X"2D",X"00",X"2B",X"60",X"93",
		X"1B",X"FF",X"73",X"A0",X"5A",X"CD",X"F3",X"75",
		X"CD",X"AC",X"4C",X"6F",X"61",X"64",X"69",X"6E",
		X"67",X"20",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"CF",X"32",X"CF",X"BD",X"CF",X"A1",X"CF",X"99",
		X"5E",X"31",X"CF",X"99",X"5E",X"30",X"CF",X"99",
		X"5E",X"29",X"CF",X"99",X"F0",X"30",X"93",X"30",
		X"1A",X"29",X"E6",X"01",X"35",X"72",X"BC",X"CF",
		X"99",X"35",X"72",X"B4",X"CF",X"99",X"5E",X"31",
		X"CF",X"99",X"5E",X"30",X"CF",X"99",X"35",X"50",
		X"E1",X"59",X"00",X"2B",X"30",X"11",X"00",X"02",
		X"2B",X"36",X"CF",X"38",X"21",X"36",X"E6",X"01",
		X"35",X"4D",X"E4",X"CF",X"5A",X"63",X"FF",X"2B",
		X"C5",X"93",X"1B",X"FF",X"74",X"A0",X"50",X"CD",
		X"C9",X"CD",X"AE",X"53",X"59",X"53",X"54",X"45",
		X"4D",X"20",X"20",X"47",X"54",X"31",X"00",X"2B",
		X"52",X"21",X"50",X"2B",X"36",X"21",X"52",X"AD",
		X"93",X"52",X"35",X"3F",X"C8",X"2B",X"C1",X"21",
		X"36",X"AD",X"93",X"36",X"FC",X"C1",X"35",X"3F",
		X"B4",X"FF",X"2B",X"C3",X"CD",X"E9",X"59",X"78",
		X"2B",X"36",X"99",X"36",X"E3",X"FE",X"2B",X"50",
		X"21",X"36",X"E3",X"07",X"F0",X"50",X"E6",X"08",
		X"35",X"4D",X"CF",X"21",X"30",X"35",X"3F",X"E4",
		X"CF",X"18",X"2B",X"C7",X"93",X"1B",X"FF",X"75",
		X"A0",X"26",X"CD",X"BF",X"75",X"93",X"56",X"11",
		X"FF",X"1F",X"F8",X"91",X"35",X"72",X"BD",X"21",
		X"CD",X"E3",X"04",X"2B",X"CD",X"F6",X"2B",X"72",
		X"21",X"CD",X"E3",X"02",X"F6",X"2B",X"74",X"CF",
		X"9B",X"63",X"FF",X"2B",X"97",X"93",X"1B",X"FF",
		X"76",X"A0",X"4B",X"CD",X"E4",X"75",X"11",X"A0",
		X"7F",X"2B",X"CD",X"CF",X"A9",X"CF",X"AB",X"21",
		X"72",X"F3",X"CD",X"93",X"CD",X"93",X"CD",X"21",
		X"74",X"F3",X"CD",X"93",X"CD",X"93",X"CD",X"11",
		X"00",X"F0",X"FA",X"74",X"E3",X"01",X"35",X"72",
		X"CA",X"59",X"07",X"FA",X"72",X"E3",X"01",X"35",
		X"3F",X"D3",X"CF",X"00",X"FD",X"04",X"68",X"18",
		X"CF",X"CF",X"AB",X"90",X"AA",X"11",X"A0",X"7F",
		X"2B",X"CD",X"F6",X"2B",X"72",X"21",X"CD",X"E3",
		X"02",X"F6",X"2B",X"74",X"63",X"FF",X"2B",X"9F",
		X"93",X"1B",X"FF",X"77",X"A0",X"5B",X"CD",X"F4",
		X"75",X"1A",X"73",X"5E",X"76",X"1A",X"74",X"5E",
		X"77",X"1A",X"75",X"2B",X"78",X"1A",X"72",X"2B",
		X"D1",X"82",X"80",X"AD",X"2B",X"72",X"59",X"00",
		X"2B",X"74",X"CF",X"7A",X"CF",X"7A",X"21",X"7C",
		X"2B",X"76",X"21",X"7E",X"2B",X"78",X"CF",X"7A",
		X"FC",X"56",X"35",X"72",X"D1",X"21",X"74",X"FC",
		X"54",X"35",X"3F",X"DE",X"21",X"72",X"2B",X"56",
		X"21",X"74",X"2B",X"54",X"CF",X"66",X"21",X"D1",
		X"82",X"7F",X"E9",X"E9",X"99",X"30",X"2B",X"D1",
		X"F6",X"2B",X"72",X"21",X"D1",X"E3",X"02",X"F6",
		X"2B",X"74",X"63",X"FF",X"2B",X"CF",X"93",X"1B",
		X"FF",X"78",X"A0",X"44",X"CD",X"B2",X"0A",X"2A",
		X"2A",X"2A",X"20",X"4D",X"65",X"6D",X"6F",X"72",
		X"79",X"20",X"63",X"61",X"72",X"64",X"0A",X"00",
		X"CF",X"32",X"59",X"00",X"5E",X"0E",X"CF",X"64",
		X"CD",X"C6",X"43",X"61",X"72",X"64",X"54",X"79",
		X"70",X"65",X"20",X"00",X"CF",X"32",X"21",X"34",
		X"CF",X"62",X"CF",X"A9",X"CF",X"6E",X"CF",X"40",
		X"35",X"72",X"D7",X"CF",X"6C",X"CF",X"89",X"CF",
		X"9D",X"35",X"72",X"E0",X"CF",X"C9",X"B4",X"80",
		X"00",X"42",X"6F",X"6F",X"74",X"00",X"00",X"00",
		X"00",X"33",X"18",X"EB",X"FB",X"EE",X"19",X"02",
		X"00",X"DD",X"21",X"11",X"35",X"56",X"0F",X"82",
		X"10",X"35",X"72",X"0F",X"11",X"45",X"E6",X"2B",
		X"24",X"B4",X"E2",X"CD",X"5F",X"21",X"30",X"E6",
		X"52",X"35",X"53",X"21",X"E3",X"32",X"2B",X"32",
		X"11",X"00",X"07",X"90",X"26",X"2B",X"32",X"11",
		X"00",X"08",X"2B",X"00",X"FD",X"04",X"68",X"18",
		X"34",X"21",X"32",X"E9",X"E9",X"99",X"32",X"99",
		X"34",X"2B",X"34",X"59",X"20",X"5E",X"24",X"21",
		X"36",X"5E",X"25",X"21",X"38",X"2B",X"28",X"E3",
		X"06",X"2B",X"38",X"11",X"E1",X"04",X"2B",X"22",
		X"59",X"FB",X"2B",X"32",X"21",X"34",X"7F",X"00",
		X"93",X"34",X"5E",X"26",X"B4",X"CB",X"93",X"28",
		X"93",X"32",X"21",X"32",X"35",X"72",X"4B",X"FF",
		X"2B",X"3A",X"CD",X"8C",X"75",X"2B",X"3C",X"21",
		X"3C",X"AD",X"35",X"3F",X"8A",X"2B",X"30",X"93",
		X"3C",X"8C",X"09",X"35",X"72",X"7D",X"21",X"38",
		X"E3",X"12",X"2B",X"38",X"90",X"66",X"8C",X"03",
		X"35",X"72",X"86",X"CF",X"3E",X"90",X"66",X"CF",
		X"3A",X"90",X"66",X"63",X"FF",X"2B",X"40",X"CD",
		X"A6",X"75",X"59",X"2D",X"2B",X"30",X"59",X"1A",
		X"2B",X"42",X"CF",X"3A",X"21",X"42",X"E6",X"01",
		X"35",X"4D",X"97",X"CF",X"3E",X"63",X"FF",X"2B",
		X"44",X"CD",X"D6",X"75",X"21",X"46",X"E6",X"06",
		X"35",X"53",X"B7",X"11",X"0B",X"20",X"90",X"BA",
		X"11",X"59",X"F0",X"2B",X"38",X"21",X"46",X"2B",
		X"42",X"11",X"00",X"08",X"99",X"38",X"2B",X"38",
		X"21",X"42",X"E6",X"01",X"35",X"53",X"BE",X"59",
		X"82",X"2B",X"30",X"CF",X"3A",X"63",X"FF",X"2B",
		X"48",X"93",X"1B",X"FF",X"03",X"00",X"A4",X"CD",
		X"9D",X"75",X"1A",X"0E",X"2B",X"36",X"CF",X"48",
		X"1A",X"11",X"8C",X"FE",X"35",X"72",X"1F",X"CF",
		X"4A",X"21",X"46",X"E6",X"05",X"35",X"4D",X"1B",
		X"E3",X"0B",X"2B",X"46",X"59",X"EF",X"5E",X"11",
		X"1A",X"11",X"8C",X"FD",X"35",X"72",X"35",X"CF",
		X"4A",X"21",X"46",X"E6",X"06",X"35",X"50",X"31",
		X"2B",X"46",X"59",X"EF",X"5E",X"11",X"1A",X"11",
		X"8C",X"FB",X"35",X"72",X"50",X"CF",X"4A",X"21",
		X"46",X"E6",X"05",X"00",X"FD",X"04",X"68",X"18",
		X"35",X"3F",X"4C",X"E6",X"06",X"35",X"3F",X"4C",
		X"93",X"46",X"59",X"EF",X"5E",X"11",X"1A",X"11",
		X"8C",X"F7",X"35",X"72",X"6D",X"CF",X"4A",X"21",
		X"46",X"35",X"3F",X"69",X"E6",X"06",X"35",X"3F",
		X"69",X"21",X"46",X"E6",X"01",X"2B",X"46",X"59",
		X"EF",X"5E",X"11",X"1A",X"11",X"82",X"80",X"35",
		X"72",X"01",X"59",X"2A",X"2B",X"36",X"CF",X"48",
		X"CD",X"94",X"0E",X"39",X"C1",X"4C",X"20",X"54",
		X"7A",X"59",X"94",X"5B",X"70",X"5A",X"F3",X"5D",
		X"38",X"85",X"19",X"98",X"8C",X"8B",X"29",X"C0",
		X"8F",X"A2",X"99",X"46",X"99",X"46",X"F6",X"2B",
		X"4C",X"63",X"FF",X"2B",X"4E",X"93",X"1B",X"FF",
		X"04",X"00",X"D6",X"CD",X"0B",X"1A",X"39",X"E3",
		X"08",X"5E",X"39",X"59",X"02",X"5E",X"38",X"FF",
		X"2B",X"3E",X"CD",X"81",X"09",X"53",X"6E",X"61",
		X"6B",X"65",X"09",X"20",X"20",X"09",X"54",X"65",
		X"74",X"72",X"6F",X"6E",X"69",X"73",X"0A",X"09",
		X"52",X"61",X"63",X"65",X"72",X"09",X"20",X"20",
		X"09",X"42",X"72",X"69",X"63",X"6B",X"73",X"0A",
		X"09",X"4D",X"61",X"6E",X"64",X"65",X"6C",X"62",
		X"72",X"6F",X"74",X"09",X"54",X"69",X"63",X"54",
		X"61",X"63",X"54",X"6F",X"65",X"0A",X"09",X"50",
		X"69",X"63",X"74",X"75",X"72",X"65",X"73",X"20",
		X"20",X"09",X"42",X"41",X"53",X"49",X"43",X"0A",
		X"09",X"43",X"72",X"65",X"64",X"69",X"74",X"73",
		X"09",X"09",X"4D",X"53",X"20",X"42",X"41",X"53",
		X"49",X"43",X"0A",X"09",X"4C",X"6F",X"61",X"64",
		X"65",X"72",X"09",X"20",X"09",X"41",X"70",X"70",
		X"6C",X"65",X"2D",X"31",X"0A",X"00",X"2B",X"50",
		X"CD",X"CF",X"55",X"73",X"65",X"20",X"5B",X"41",
		X"72",X"72",X"6F",X"77",X"73",X"5D",X"20",X"74",
		X"6F",X"20",X"73",X"00",X"FD",X"04",X"68",X"18",
		X"65",X"6C",X"65",X"63",X"74",X"0A",X"50",X"72",
		X"65",X"73",X"73",X"20",X"5B",X"41",X"5D",X"20",
		X"74",X"6F",X"20",X"73",X"74",X"61",X"72",X"74",
		X"20",X"70",X"72",X"6F",X"67",X"72",X"61",X"6D",
		X"0A",X"0A",X"48",X"6F",X"6C",X"64",X"20",X"5B",
		X"53",X"74",X"61",X"72",X"74",X"5D",X"20",X"66",
		X"6F",X"72",X"20",X"72",X"65",X"73",X"65",X"74",
		X"00",X"2B",X"52",X"93",X"1B",X"FF",X"05",X"00",
		X"B7",X"CD",X"11",X"75",X"21",X"38",X"E6",X"0C",
		X"2B",X"38",X"59",X"20",X"2B",X"30",X"CF",X"3A",
		X"CF",X"3A",X"63",X"FF",X"2B",X"4A",X"CD",X"30",
		X"75",X"59",X"2A",X"2B",X"36",X"CF",X"44",X"59",
		X"0F",X"2B",X"36",X"21",X"50",X"CF",X"40",X"59",
		X"2A",X"2B",X"36",X"CF",X"44",X"21",X"52",X"CF",
		X"40",X"63",X"FF",X"2B",X"54",X"1A",X"21",X"88",
		X"03",X"5E",X"21",X"59",X"5A",X"5E",X"2C",X"11",
		X"02",X"20",X"2B",X"38",X"CF",X"54",X"59",X"00",
		X"2B",X"46",X"CF",X"4E",X"11",X"00",X"08",X"2B",
		X"28",X"11",X"01",X"88",X"2B",X"32",X"11",X"80",
		X"FF",X"2B",X"42",X"21",X"38",X"E3",X"30",X"F8",
		X"42",X"2B",X"56",X"11",X"E1",X"04",X"2B",X"22",
		X"59",X"20",X"5E",X"24",X"5E",X"25",X"21",X"28",
		X"E3",X"30",X"F8",X"42",X"FC",X"56",X"35",X"3F",
		X"7F",X"1A",X"59",X"8C",X"78",X"35",X"3F",X"7F",
		X"B4",X"CB",X"11",X"00",X"08",X"99",X"28",X"2B",
		X"28",X"35",X"4D",X"6D",X"99",X"32",X"2B",X"28",
		X"82",X"FF",X"8C",X"A0",X"35",X"72",X"6B",X"59",
		X"AD",X"2B",X"22",X"21",X"4C",X"2B",X"24",X"11",
		X"00",X"02",X"2B",X"1A",X"21",X"46",X"E6",X"0A",
		X"35",X"3F",X"AA",X"E6",X"01",X"35",X"72",X"B3",
		X"1A",X"21",X"82",X"F8",X"5E",X"21",X"B4",X"E2",
		X"00",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"4D",X"61",X"69",X"6E",X"00",X"00",X"00",X"00",
		X"CF",X"18",X"F5",X"FB",X"EE",X"19",X"02",X"00",
		X"F3",X"11",X"F8",X"01",X"2B",X"30",X"CD",X"75",
		X"75",X"1A",X"01",X"E6",X"01",X"82",X"FF",X"E3",
		X"01",X"2B",X"32",X"11",X"09",X"0B",X"2B",X"22",
		X"59",X"AA",X"5E",X"7C",X"59",X"7C",X"B4",X"FA",
		X"1A",X"7C",X"8C",X"AA",X"35",X"3F",X"2A",X"59",
		X"00",X"F0",X"30",X"90",X"54",X"11",X"24",X"80",
		X"2B",X"34",X"59",X"BC",X"B4",X"FA",X"21",X"34",
		X"AD",X"8C",X"FF",X"F0",X"34",X"2B",X"24",X"8C",
		X"FF",X"F0",X"34",X"FC",X"24",X"35",X"3F",X"4F",
		X"59",X"31",X"2B",X"36",X"CF",X"38",X"59",X"70",
		X"2B",X"32",X"11",X"7C",X"80",X"B4",X"FA",X"11",
		X"2F",X"2F",X"2B",X"36",X"21",X"32",X"93",X"36",
		X"E6",X"28",X"35",X"53",X"5B",X"E3",X"28",X"93",
		X"37",X"E6",X"04",X"35",X"53",X"64",X"CF",X"38",
		X"1A",X"37",X"2B",X"36",X"CF",X"38",X"63",X"FF",
		X"2B",X"3A",X"CD",X"9D",X"75",X"2B",X"3C",X"21",
		X"3C",X"AD",X"35",X"3F",X"9B",X"2B",X"36",X"8C",
		X"0A",X"35",X"3F",X"8D",X"CF",X"38",X"90",X"97",
		X"59",X"02",X"5E",X"3E",X"1A",X"3F",X"E3",X"08",
		X"5E",X"3F",X"93",X"3C",X"90",X"7C",X"63",X"FF",
		X"2B",X"40",X"CD",X"EC",X"1A",X"36",X"E6",X"52",
		X"35",X"53",X"B1",X"E3",X"32",X"2B",X"32",X"11",
		X"00",X"07",X"90",X"B6",X"2B",X"32",X"11",X"00",
		X"08",X"2B",X"42",X"21",X"32",X"E9",X"E9",X"99",
		X"32",X"99",X"42",X"2B",X"42",X"11",X"E1",X"04",
		X"2B",X"22",X"11",X"20",X"3F",X"2B",X"24",X"21",
		X"3E",X"2B",X"28",X"E3",X"06",X"2B",X"3E",X"59",
		X"05",X"2B",X"32",X"21",X"42",X"7F",X"00",X"5E",
		X"26",X"B4",X"CB",X"93",X"42",X"93",X"28",X"21",
		X"32",X"E6",X"01",X"00",X"FD",X"04",X"68",X"18",
		X"35",X"4D",X"D6",X"FF",X"2B",X"38",X"93",X"1B",
		X"FF",X"03",X"00",X"EA",X"CD",X"37",X"2B",X"32",
		X"88",X"FF",X"8C",X"FF",X"88",X"FA",X"2B",X"44",
		X"1A",X"32",X"2B",X"32",X"59",X"00",X"F0",X"44",
		X"93",X"44",X"59",X"03",X"F0",X"44",X"93",X"44",
		X"11",X"00",X"09",X"99",X"32",X"7F",X"00",X"F0",
		X"44",X"93",X"44",X"11",X"00",X"09",X"99",X"32",
		X"7F",X"01",X"F0",X"44",X"93",X"44",X"F0",X"44",
		X"93",X"44",X"F0",X"44",X"FF",X"2B",X"46",X"CD",
		X"C9",X"75",X"59",X"10",X"2B",X"42",X"59",X"0A",
		X"2B",X"32",X"CF",X"48",X"21",X"32",X"E6",X"01",
		X"35",X"4D",X"42",X"11",X"09",X"0B",X"2B",X"22",
		X"11",X"78",X"80",X"B4",X"FA",X"CD",X"61",X"FF",
		X"FF",X"40",X"00",X"00",X"00",X"00",X"95",X"2B",
		X"44",X"59",X"81",X"2B",X"34",X"59",X"08",X"2B",
		X"32",X"21",X"44",X"AD",X"93",X"44",X"F0",X"34",
		X"93",X"34",X"21",X"32",X"E6",X"01",X"35",X"4D",
		X"69",X"59",X"81",X"2B",X"24",X"E3",X"08",X"2B",
		X"26",X"11",X"15",X"0B",X"2B",X"22",X"B4",X"CB",
		X"59",X"10",X"2B",X"32",X"CF",X"48",X"82",X"80",
		X"35",X"3F",X"9C",X"21",X"32",X"E6",X"01",X"35",
		X"4D",X"8C",X"11",X"09",X"0B",X"2B",X"22",X"11",
		X"7C",X"80",X"B4",X"FA",X"1A",X"2A",X"35",X"3F",
		X"C7",X"8C",X"01",X"35",X"72",X"C0",X"11",X"33",
		X"EB",X"2B",X"24",X"11",X"00",X"02",X"2B",X"1A",
		X"59",X"AD",X"2B",X"22",X"B4",X"E2",X"21",X"42",
		X"E6",X"01",X"35",X"4D",X"3E",X"63",X"FF",X"2B",
		X"4A",X"CD",X"E3",X"59",X"FF",X"5E",X"2A",X"59",
		X"2A",X"2B",X"24",X"E3",X"01",X"2B",X"26",X"11",
		X"15",X"0B",X"2B",X"22",X"B4",X"CB",X"1A",X"2A",
		X"FF",X"2B",X"48",X"93",X"1B",X"FF",X"04",X"00",
		X"D6",X"11",X"0F",X"00",X"FD",X"04",X"68",X"18",
		X"0B",X"2B",X"22",X"59",X"00",X"B4",X"F5",X"11",
		X"12",X"0B",X"2B",X"22",X"59",X"00",X"B4",X"F7",
		X"B4",X"F7",X"B4",X"F7",X"B4",X"F7",X"11",X"58",
		X"01",X"CF",X"46",X"11",X"70",X"02",X"CF",X"46",
		X"11",X"78",X"03",X"CF",X"46",X"11",X"7E",X"04",
		X"CF",X"46",X"11",X"00",X"01",X"2B",X"44",X"11",
		X"00",X"08",X"2B",X"34",X"1A",X"35",X"F0",X"44",
		X"93",X"44",X"59",X"00",X"F0",X"44",X"93",X"44",
		X"93",X"35",X"21",X"34",X"35",X"4D",X"34",X"11",
		X"03",X"0B",X"2B",X"22",X"59",X"20",X"5E",X"25",
		X"11",X"00",X"08",X"2B",X"44",X"2B",X"26",X"59",
		X"A0",X"5E",X"24",X"B4",X"F3",X"11",X"00",X"01",
		X"99",X"44",X"35",X"4D",X"53",X"1A",X"2E",X"82",
		X"80",X"35",X"72",X"70",X"5E",X"2E",X"5E",X"2D",
		X"59",X"09",X"5E",X"2F",X"11",X"14",X"08",X"2B",
		X"3E",X"CD",X"89",X"2A",X"2A",X"2A",X"20",X"47",
		X"69",X"67",X"61",X"74",X"72",X"6F",X"6E",X"20",
		X"00",X"CF",X"40",X"CF",X"3A",X"CD",X"B1",X"4B",
		X"20",X"2A",X"2A",X"2A",X"20",X"0A",X"20",X"54",
		X"54",X"4C",X"20",X"6D",X"69",X"63",X"72",X"6F",
		X"63",X"6F",X"6D",X"70",X"75",X"74",X"65",X"72",
		X"20",X"52",X"4F",X"4D",X"20",X"76",X"35",X"61",
		X"00",X"CF",X"40",X"11",X"00",X"0B",X"2B",X"22",
		X"59",X"01",X"B4",X"E6",X"21",X"30",X"AD",X"35",
		X"3F",X"C4",X"CF",X"4A",X"11",X"CF",X"F5",X"2B",
		X"24",X"11",X"00",X"02",X"2B",X"1A",X"59",X"AD",
		X"2B",X"22",X"B4",X"E2",X"00",X"DB",X"24",X"00",
		X"18",X"0E",X"00",X"00",X"E0",X"FB",X"00",X"00",
		X"52",X"65",X"73",X"65",X"74",X"00",X"00",X"00",
		X"0E",X"18",X"F9",X"FB",X"EE",X"19",X"03",X"CB",
		X"EA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FD",X"04",X"68",X"18",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		X"69",X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",
		X"21",X"69",X"61",X"72",X"6E",X"47",X"67",X"74",
		X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",X"67",
		X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",X"47",
		X"67",X"74",X"6F",X"21",X"69",X"61",X"72",X"6E",
		X"47",X"67",X"74",X"6F",X"21",X"69",X"61",X"72",
		X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",X"61",
		X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",X"69",
		X"61",X"72",X"6E",X"47",X"67",X"74",X"6F",X"21",
		others => (others => '0'));
	signal q0_reg : rom_data_elem_t;
	signal q1_reg : rom_data_elem_t;
begin
	q(7 downto 0) <= q0_reg;
	q(15 downto 8) <= q1_reg;
	process(a)
	begin
		q0_reg <= rom_data_byte0(to_integer(a));
		q1_reg <= rom_data_byte1(to_integer(a));
	end process;
end architecture;
